-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.43919902411519324]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_d7300028 is
port(
 clk : in std_logic;
 elem_val : in unsigned(31 downto 0);
 ref_toks_0 : in chacha20_state;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint32_t_array_16_t);
end VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_d7300028;
architecture arch of VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_d7300028 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 1;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue : unsigned(31 downto 0);
signal REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue : unsigned(31 downto 0);
signal COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse : unsigned(31 downto 0);
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint32_t_array_16_t is
 
  variable base : uint32_t_array_16_t; 
  variable return_output : uint32_t_array_16_t;
begin
      base.data(0) := ref_toks_0;
      base.data(3) := ref_toks_1;
      base.data(9) := ref_toks_2;
      base.data(6) := ref_toks_3;
      base.data(12) := ref_toks_4;
      base.data(15) := ref_toks_5;
      base.data(4) := ref_toks_6;
      base.data(1) := ref_toks_7;
      base.data(7) := ref_toks_8;
      base.data(10) := ref_toks_9;
      base.data(13) := ref_toks_10;
      base.data(2) := ref_toks_11;
      base.data(5) := ref_toks_12;
      base.data(11) := ref_toks_13;
      base.data(8) := ref_toks_14;
      base.data(14) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d : 1 clocks latency
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_d4eec02f port map (
clk,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413 : entity work.BIN_OP_EQ_uint4_t_uint2_t_1CLK_ef275fc6 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5 : 0 clocks latency
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c : 0 clocks latency
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140 : entity work.BIN_OP_EQ_uint4_t_uint3_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd : 0 clocks latency
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e : 0 clocks latency
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877 : 0 clocks latency
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971 : entity work.BIN_OP_EQ_uint4_t_uint3_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78 : 0 clocks latency
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2 : 1 clocks latency
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_d4eec02f port map (
clk,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75 : entity work.BIN_OP_EQ_uint4_t_uint3_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b : 0 clocks latency
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc : 0 clocks latency
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53 : 0 clocks latency
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793 : entity work.BIN_OP_EQ_uint4_t_uint2_t_1CLK_ef275fc6 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845 : 0 clocks latency
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555 : entity work.BIN_OP_EQ_uint4_t_uint3_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee : 0 clocks latency
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51 : 0 clocks latency
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c : 0 clocks latency
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92 : 1 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92 : entity work.BIN_OP_EQ_uint4_t_uint4_t_1CLK_fdcb26f0 port map (
clk,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102 : 0 clocks latency
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- Registers
 -- Stage 0
 REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue,
 REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse,
 REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue,
 REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse,
 REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue,
 REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse,
 REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue,
 REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse,
 REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue,
 REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse,
 REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue,
 REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse,
 REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue,
 REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse,
 REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue,
 REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse,
 REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue,
 REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse,
 REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue,
 REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse,
 REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue,
 REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse,
 REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue,
 REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse,
 REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue,
 REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse,
 REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue,
 REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(31 downto 0);
 variable VAR_ref_toks_0 : chacha20_state;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint32_t_array_16_t;
 variable VAR_base : chacha20_state;
 variable VAR_rv : uint32_t_array_16_t;
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5144_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_ac05_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_ecef_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b9bf_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_0298_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c16_2e43_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_afa7_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_e8b5_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_4546_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_3ca4_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_097f_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_890d_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_2aa8_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c16_ba98_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_adc6_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_7b50_return_output : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_2a86_return_output : uint32_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right := to_unsigned(14, 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left := VAR_var_dim_0;
     -- CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5144] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5144_return_output := VAR_ref_toks_0.state(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_097f] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_097f_return_output := VAR_ref_toks_0.state(13);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_afa7] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_afa7_return_output := VAR_ref_toks_0.state(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_ac05] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_ac05_return_output := VAR_ref_toks_0.state(3);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_4546] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_4546_return_output := VAR_ref_toks_0.state(7);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_7b50] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_7b50_return_output := VAR_ref_toks_0.state(14);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b9bf] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b9bf_return_output := VAR_ref_toks_0.state(6);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_adc6] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_adc6_return_output := VAR_ref_toks_0.state(8);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_ecef] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_ecef_return_output := VAR_ref_toks_0.state(9);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c16_ba98] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c16_ba98_return_output := VAR_ref_toks_0.state(11);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_890d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_890d_return_output := VAR_ref_toks_0.state(2);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_2aa8] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_2aa8_return_output := VAR_ref_toks_0.state(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_right;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c16_2e43] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c16_2e43_return_output := VAR_ref_toks_0.state(15);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9] LATENCY=1
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_right;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_3ca4] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_3ca4_return_output := VAR_ref_toks_0.state(10);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_0298] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_0298_return_output := VAR_ref_toks_0.state(12);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_e8b5] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_e8b5_return_output := VAR_ref_toks_0.state(1);

     -- Submodule level 1
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_ac79_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_ef2c_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5144_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_3ca4_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c16_ba98_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_0298_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_097f_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_7b50_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c16_2e43_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_e8b5_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_890d_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_ac05_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_afa7_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_2aa8_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b9bf_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_4546_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c15_adc6_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c15_ecef_return_output;
     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2] LATENCY=1
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_iffalse;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d] LATENCY=1
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_iffalse;

     -- Write to comb signals
     COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue;
     COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse;
     COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue;
     COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse;
     COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue;
     COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse;
     COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue;
     COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse;
     COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue;
     COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse;
     COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue;
     COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse;
     COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue;
     COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse;
     COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue;
     COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse;
     COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue;
     COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse;
     COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue;
     COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse;
     COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue;
     COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse;
     COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue;
     COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse;
     COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue;
     COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse;
     COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue;
     COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue := REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse := REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue := REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse := REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue := REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse := REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue := REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse := REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue := REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse := REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue := REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse := REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue := REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse := REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue := REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse := REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue := REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse := REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue := REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse := REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue := REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse := REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue := REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse := REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue := REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse := REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue := REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse := REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse;
     -- Submodule outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output;

     -- Submodule level 0
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_b793_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_b555_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_c813_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_00f9_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6e92_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_3413_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_ffb8_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_9140_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_f83e_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_8ab8_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_e971_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_bd75_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_fcc2_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_4c64_return_output;
     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_2a86] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_2a86_return_output := CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0(
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_828d_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_35b2_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_return_output);

     -- Submodule level 2
     VAR_return_output := VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_53b0_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_2a86_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue <= COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iftrue;
     REG_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse <= COMB_STAGE0_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_2be5_iffalse;
     REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue <= COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iftrue;
     REG_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse <= COMB_STAGE0_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_1c0c_iffalse;
     REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue <= COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iftrue;
     REG_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse <= COMB_STAGE0_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_0bfd_iffalse;
     REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue <= COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iftrue;
     REG_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse <= COMB_STAGE0_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_801e_iffalse;
     REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue <= COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iftrue;
     REG_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse <= COMB_STAGE0_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_7877_iffalse;
     REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue <= COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iftrue;
     REG_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse <= COMB_STAGE0_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_0b78_iffalse;
     REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue <= COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iftrue;
     REG_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse <= COMB_STAGE0_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_f80b_iffalse;
     REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue <= COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iftrue;
     REG_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse <= COMB_STAGE0_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_ecfc_iffalse;
     REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue <= COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iftrue;
     REG_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse <= COMB_STAGE0_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_4d53_iffalse;
     REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue <= COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iftrue;
     REG_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse <= COMB_STAGE0_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_c845_iffalse;
     REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue <= COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iftrue;
     REG_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse <= COMB_STAGE0_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_a0ee_iffalse;
     REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue <= COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iftrue;
     REG_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse <= COMB_STAGE0_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_cc51_iffalse;
     REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue <= COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iftrue;
     REG_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse <= COMB_STAGE0_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_664c_iffalse;
     REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue <= COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iftrue;
     REG_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse <= COMB_STAGE0_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_2102_iffalse;
 end if;
end process;

end arch;
