module imem (
	clk,
	arst_n,
	rvld,
	rrdy,
	raddr,
	rdat,
	we,
	waddr,
	wdat
);
	parameter signed [31:0] NUM_WORDS = 8192;
	input wire clk;
	input wire arst_n;
	input wire rvld;
	output reg rrdy;
	input wire [31:2] raddr;
	output reg [31:0] rdat;
	input wire we;
	input wire [31:2] waddr;
	input wire [31:0] wdat;
	localparam ADDR_MSB = $clog2(NUM_WORDS) + 1;
	reg [31:0] mem [0:NUM_WORDS - 1];
	wire [ADDR_MSB:2] raddr_int;
	wire [ADDR_MSB:2] waddr_int;
	assign raddr_int = raddr[ADDR_MSB:2];
	assign waddr_int = waddr[ADDR_MSB:2];
	initial begin
		mem['h0] = 32'h00001517;
		mem['h1] = 32'h23050513;
		mem['h2] = 32'h10000597;
		mem['h3] = 32'hff858593;
		mem['h4] = 32'h10000617;
		mem['h5] = 32'h00860613;
		mem['h6] = 32'h00c5dc63;
		mem['h7] = 32'h00052683;
		mem['h8] = 32'h00d5a023;
		mem['h9] = 32'h00450513;
		mem['ha] = 32'h00458593;
		mem['hb] = 32'hfec5c8e3;
		mem['hc] = 32'h10000517;
		mem['hd] = 32'hfe850513;
		mem['he] = 32'h10001597;
		mem['hf] = 32'h3f458593;
		mem['h10] = 32'h00b55863;
		mem['h11] = 32'h00052023;
		mem['h12] = 32'h00450513;
		mem['h13] = 32'hfeb54ce3;
		mem['h14] = 32'h10008117;
		mem['h15] = 32'hfb010113;
		mem['h16] = 32'h10000197;
		mem['h17] = 32'h7c018193;
		mem['h18] = 32'h00a54533;
		mem['h19] = 32'h00b5c5b3;
		mem['h1a] = 32'h00c64633;
		mem['h1b] = 32'h530000ef;
		mem['h1c] = 32'h0000006f;
		mem['h1d] = 32'h00452783;
		mem['h1e] = 32'h0087a783;
		mem['h1f] = 32'h0007a783;
		mem['h20] = 32'h0007a783;
		mem['h21] = 32'hfe07c8e3;
		mem['h22] = 32'h00452783;
		mem['h23] = 32'h0087a783;
		mem['h24] = 32'h0007a783;
		mem['h25] = 32'h00b78023;
		mem['h26] = 32'h00008067;
		mem['h27] = 32'h0a058a63;
		mem['h28] = 32'hfe010113;
		mem['h29] = 32'h00912a23;
		mem['h2a] = 32'h00058493;
		mem['h2b] = 32'h01212823;
		mem['h2c] = 32'h00a00593;
		mem['h2d] = 32'h00050913;
		mem['h2e] = 32'h00048513;
		mem['h2f] = 32'h00812c23;
		mem['h30] = 32'h00112e23;
		mem['h31] = 32'h01312623;
		mem['h32] = 32'h01412423;
		mem['h33] = 32'h701000ef;
		mem['h34] = 32'h01051513;
		mem['h35] = 32'h01055513;
		mem['h36] = 32'h00100413;
		mem['h37] = 32'h06857e63;
		mem['h38] = 32'h00900a13;
		mem['h39] = 32'h00040593;
		mem['h3a] = 32'h00048513;
		mem['h3b] = 32'h6e1000ef;
		mem['h3c] = 32'h03050593;
		mem['h3d] = 32'h0ff5f593;
		mem['h3e] = 32'h00090513;
		mem['h3f] = 32'hf79ff0ef;
		mem['h40] = 32'h00040593;
		mem['h41] = 32'h00048513;
		mem['h42] = 32'h70d000ef;
		mem['h43] = 32'h01051493;
		mem['h44] = 32'h00a00593;
		mem['h45] = 32'h00040513;
		mem['h46] = 32'h6b5000ef;
		mem['h47] = 32'h00040993;
		mem['h48] = 32'h01051413;
		mem['h49] = 32'h0104d493;
		mem['h4a] = 32'h01045413;
		mem['h4b] = 32'hfb3a6ce3;
		mem['h4c] = 32'h01c12083;
		mem['h4d] = 32'h01812403;
		mem['h4e] = 32'h01412483;
		mem['h4f] = 32'h01012903;
		mem['h50] = 32'h00c12983;
		mem['h51] = 32'h00812a03;
		mem['h52] = 32'h02010113;
		mem['h53] = 32'h00008067;
		mem['h54] = 32'h03000593;
		mem['h55] = 32'hf21ff06f;
		mem['h56] = 32'h00241793;
		mem['h57] = 32'h00f40433;
		mem['h58] = 32'h00141413;
		mem['h59] = 32'h01041413;
		mem['h5a] = 32'h01045413;
		mem['h5b] = 32'hf71ff06f;
		mem['h5c] = 32'hff010113;
		mem['h5d] = 32'h00812423;
		mem['h5e] = 32'h00912223;
		mem['h5f] = 32'h00112623;
		mem['h60] = 32'h00050493;
		mem['h61] = 32'h00058413;
		mem['h62] = 32'h00044583;
		mem['h63] = 32'h00058a63;
		mem['h64] = 32'h00048513;
		mem['h65] = 32'h00140413;
		mem['h66] = 32'heddff0ef;
		mem['h67] = 32'hfedff06f;
		mem['h68] = 32'h00c12083;
		mem['h69] = 32'h00812403;
		mem['h6a] = 32'h00412483;
		mem['h6b] = 32'h01010113;
		mem['h6c] = 32'h00008067;
		mem['h6d] = 32'hff010113;
		mem['h6e] = 32'h00112623;
		mem['h6f] = 32'h00812423;
		mem['h70] = 32'h00912223;
		mem['h71] = 32'h00058493;
		mem['h72] = 32'h0005c583;
		mem['h73] = 32'h00050413;
		mem['h74] = 32'hecdff0ef;
		mem['h75] = 32'h00040513;
		mem['h76] = 32'h02e00593;
		mem['h77] = 32'he99ff0ef;
		mem['h78] = 32'h0014c583;
		mem['h79] = 32'h00040513;
		mem['h7a] = 32'heb5ff0ef;
		mem['h7b] = 32'h00040513;
		mem['h7c] = 32'h02e00593;
		mem['h7d] = 32'he81ff0ef;
		mem['h7e] = 32'h0024c583;
		mem['h7f] = 32'h00040513;
		mem['h80] = 32'he9dff0ef;
		mem['h81] = 32'h00040513;
		mem['h82] = 32'h02e00593;
		mem['h83] = 32'he69ff0ef;
		mem['h84] = 32'h00040513;
		mem['h85] = 32'h00812403;
		mem['h86] = 32'h0034c583;
		mem['h87] = 32'h00c12083;
		mem['h88] = 32'h00412483;
		mem['h89] = 32'h01010113;
		mem['h8a] = 32'he75ff06f;
		mem['h8b] = 32'h00100613;
		mem['h8c] = 32'h00010837;
		mem['h8d] = 32'h00050713;
		mem['h8e] = 32'h00000793;
		mem['h8f] = 32'h40a60633;
		mem['h90] = 32'hfff80893;
		mem['h91] = 32'h00e606b3;
		mem['h92] = 32'h02b6f663;
		mem['h93] = 32'h00074683;
		mem['h94] = 32'h00174303;
		mem['h95] = 32'h00869693;
		mem['h96] = 32'h0066e6b3;
		mem['h97] = 32'h00d787b3;
		mem['h98] = 32'h0107e663;
		mem['h99] = 32'h0117f7b3;
		mem['h9a] = 32'h00178793;
		mem['h9b] = 32'h00270713;
		mem['h9c] = 32'hfd5ff06f;
		mem['h9d] = 32'hffe5f713;
		mem['h9e] = 32'h02b77463;
		mem['h9f] = 32'h00e50533;
		mem['ha0] = 32'h00054703;
		mem['ha1] = 32'h00871713;
		mem['ha2] = 32'h00e787b3;
		mem['ha3] = 32'h00010737;
		mem['ha4] = 32'h00e7e863;
		mem['ha5] = 32'h01079793;
		mem['ha6] = 32'h0107d793;
		mem['ha7] = 32'h00178793;
		mem['ha8] = 32'hfff7c513;
		mem['ha9] = 32'h01051513;
		mem['haa] = 32'h01055513;
		mem['hab] = 32'h00008067;
		mem['hac] = 32'h100016b7;
		mem['had] = 32'h4286a703;
		mem['hae] = 32'h100017b7;
		mem['haf] = 32'hc2878793;
		mem['hb0] = 32'h00f707b3;
		mem['hb1] = 32'h00a70733;
		mem['hb2] = 32'h42e6a423;
		mem['hb3] = 32'h000016b7;
		mem['hb4] = 32'h80068693;
		mem['hb5] = 32'h00e6d463;
		mem['hb6] = 32'h00100073;
		mem['hb7] = 32'h00078513;
		mem['hb8] = 32'h00008067;
		mem['hb9] = 32'hff010113;
		mem['hba] = 32'h00812423;
		mem['hbb] = 32'h00001437;
		mem['hbc] = 32'h07840413;
		mem['hbd] = 32'h0045d793;
		mem['hbe] = 32'h00f407b3;
		mem['hbf] = 32'h00912223;
		mem['hc0] = 32'h00058493;
		mem['hc1] = 32'h0007c583;
		mem['hc2] = 32'h00f4f493;
		mem['hc3] = 32'h01212023;
		mem['hc4] = 32'h00112623;
		mem['hc5] = 32'h00050913;
		mem['hc6] = 32'h00940433;
		mem['hc7] = 32'hd59ff0ef;
		mem['hc8] = 32'h00044583;
		mem['hc9] = 32'h00812403;
		mem['hca] = 32'h00c12083;
		mem['hcb] = 32'h00412483;
		mem['hcc] = 32'h00090513;
		mem['hcd] = 32'h00012903;
		mem['hce] = 32'h01010113;
		mem['hcf] = 32'hd39ff06f;
		mem['hd0] = 32'h00052783;
		mem['hd1] = 32'h0007a783;
		mem['hd2] = 32'h0187a783;
		mem['hd3] = 32'h0007a783;
		mem['hd4] = 32'h0007a783;
		mem['hd5] = 32'h0017f793;
		mem['hd6] = 32'h1e078e63;
		mem['hd7] = 32'h00052783;
		mem['hd8] = 32'hffff8637;
		mem['hd9] = 32'hffff08b7;
		mem['hda] = 32'h0007a783;
		mem['hdb] = 32'hfff60613;
		mem['hdc] = 32'h0107a783;
		mem['hdd] = 32'h0007a683;
		mem['hde] = 32'h0005c783;
		mem['hdf] = 32'h0077f713;
		mem['he0] = 32'h0006a783;
		mem['he1] = 32'hff87f793;
		mem['he2] = 32'h00e7e7b3;
		mem['he3] = 32'h00f6a023;
		mem['he4] = 32'h00052783;
		mem['he5] = 32'h0007a783;
		mem['he6] = 32'h0107a783;
		mem['he7] = 32'h0007a683;
		mem['he8] = 32'h0015c783;
		mem['he9] = 32'h0077f793;
		mem['hea] = 32'h00379713;
		mem['heb] = 32'h0006a783;
		mem['hec] = 32'hfc77f793;
		mem['hed] = 32'h00e7e7b3;
		mem['hee] = 32'h00f6a023;
		mem['hef] = 32'h00052783;
		mem['hf0] = 32'h0007a783;
		mem['hf1] = 32'h0107a783;
		mem['hf2] = 32'h0007a683;
		mem['hf3] = 32'h0025c783;
		mem['hf4] = 32'h0017f793;
		mem['hf5] = 32'h00679713;
		mem['hf6] = 32'h0006a783;
		mem['hf7] = 32'hfbf7f793;
		mem['hf8] = 32'h00e7e7b3;
		mem['hf9] = 32'h00f6a023;
		mem['hfa] = 32'h00052783;
		mem['hfb] = 32'h0007a783;
		mem['hfc] = 32'h0107a783;
		mem['hfd] = 32'h0007a683;
		mem['hfe] = 32'h0035c783;
		mem['hff] = 32'h0017f793;
		mem['h100] = 32'h00779713;
		mem['h101] = 32'h0006a783;
		mem['h102] = 32'hf7f7f793;
		mem['h103] = 32'h00e7e7b3;
		mem['h104] = 32'h00f6a023;
		mem['h105] = 32'h00858713;
		mem['h106] = 32'h00000793;
		mem['h107] = 32'h00052683;
		mem['h108] = 32'h00072803;
		mem['h109] = 32'h01078793;
		mem['h10a] = 32'h0006a683;
		mem['h10b] = 32'h01070713;
		mem['h10c] = 32'h0006a683;
		mem['h10d] = 32'h0006a683;
		mem['h10e] = 32'h0106a023;
		mem['h10f] = 32'h00052683;
		mem['h110] = 32'hff472803;
		mem['h111] = 32'h0006a683;
		mem['h112] = 32'h0046a683;
		mem['h113] = 32'h0006a683;
		mem['h114] = 32'h0106a023;
		mem['h115] = 32'h00052683;
		mem['h116] = 32'hff872803;
		mem['h117] = 32'h0006a683;
		mem['h118] = 32'h0086a683;
		mem['h119] = 32'h0006a683;
		mem['h11a] = 32'h0106a023;
		mem['h11b] = 32'h00052683;
		mem['h11c] = 32'hffc72803;
		mem['h11d] = 32'h0006a683;
		mem['h11e] = 32'h00c6a683;
		mem['h11f] = 32'h0006a683;
		mem['h120] = 32'h0106a023;
		mem['h121] = 32'h0045a683;
		mem['h122] = 32'h04d7fe63;
		mem['h123] = 32'h00052683;
		mem['h124] = 32'h0006a683;
		mem['h125] = 32'h0106a683;
		mem['h126] = 32'h0006a803;
		mem['h127] = 32'h00082683;
		mem['h128] = 32'h0116e6b3;
		mem['h129] = 32'h00d82023;
		mem['h12a] = 32'h00052683;
		mem['h12b] = 32'h0006a683;
		mem['h12c] = 32'h0106a683;
		mem['h12d] = 32'h0006a803;
		mem['h12e] = 32'h00082683;
		mem['h12f] = 32'h00c6f6b3;
		mem['h130] = 32'h00d82023;
		mem['h131] = 32'h00052683;
		mem['h132] = 32'h0006a683;
		mem['h133] = 32'h0146a683;
		mem['h134] = 32'h0006a803;
		mem['h135] = 32'h00082683;
		mem['h136] = 32'h0016e693;
		mem['h137] = 32'h00d82023;
		mem['h138] = 32'hf3dff06f;
		mem['h139] = 32'h00052703;
		mem['h13a] = 32'h40d787b3;
		mem['h13b] = 32'h00072703;
		mem['h13c] = 32'h01072703;
		mem['h13d] = 32'h00072603;
		mem['h13e] = 32'h00010737;
		mem['h13f] = 32'hfff70693;
		mem['h140] = 32'h00062703;
		mem['h141] = 32'h40f6d7b3;
		mem['h142] = 32'h01079793;
		mem['h143] = 32'h00d77733;
		mem['h144] = 32'h00f767b3;
		mem['h145] = 32'h00f62023;
		mem['h146] = 32'h00052783;
		mem['h147] = 32'h000086b7;
		mem['h148] = 32'h0007a783;
		mem['h149] = 32'h0107a783;
		mem['h14a] = 32'h0007a703;
		mem['h14b] = 32'h00072783;
		mem['h14c] = 32'h00d7e7b3;
		mem['h14d] = 32'h00f72023;
		mem['h14e] = 32'h00052783;
		mem['h14f] = 32'h0007a783;
		mem['h150] = 32'h0147a783;
		mem['h151] = 32'h0007a703;
		mem['h152] = 32'h00072783;
		mem['h153] = 32'h0017e793;
		mem['h154] = 32'h00f72023;
		mem['h155] = 32'h00008067;
		mem['h156] = 32'h0ff5f593;
		mem['h157] = 32'h00000793;
		mem['h158] = 32'h00c78a63;
		mem['h159] = 32'h00f50733;
		mem['h15a] = 32'h00b70023;
		mem['h15b] = 32'h00178793;
		mem['h15c] = 32'hff1ff06f;
		mem['h15d] = 32'h00008067;
		mem['h15e] = 32'h00000793;
		mem['h15f] = 32'h00c78e63;
		mem['h160] = 32'h00f58733;
		mem['h161] = 32'h00074683;
		mem['h162] = 32'h00f50733;
		mem['h163] = 32'h00178793;
		mem['h164] = 32'h00d70023;
		mem['h165] = 32'hfe9ff06f;
		mem['h166] = 32'h00008067;
		mem['h167] = 32'hf9010113;
		mem['h168] = 32'h02800513;
		mem['h169] = 32'h06112623;
		mem['h16a] = 32'h06812423;
		mem['h16b] = 32'h06912223;
		mem['h16c] = 32'h07212023;
		mem['h16d] = 32'h05312e23;
		mem['h16e] = 32'h05412c23;
		mem['h16f] = 32'h05512a23;
		mem['h170] = 32'h05612823;
		mem['h171] = 32'h05712623;
		mem['h172] = 32'h05812423;
		mem['h173] = 32'h05912223;
		mem['h174] = 32'h05a12023;
		mem['h175] = 32'h03b12e23;
		mem['h176] = 32'hcd9ff0ef;
		mem['h177] = 32'h00050413;
		mem['h178] = 32'h00800513;
		mem['h179] = 32'hccdff0ef;
		mem['h17a] = 32'h00050993;
		mem['h17b] = 32'h01c00513;
		mem['h17c] = 32'hcc1ff0ef;
		mem['h17d] = 32'h00050913;
		mem['h17e] = 32'h00400513;
		mem['h17f] = 32'h200004b7;
		mem['h180] = 32'hcb1ff0ef;
		mem['h181] = 32'h00952023;
		mem['h182] = 32'h00a92023;
		mem['h183] = 32'h00400513;
		mem['h184] = 32'hca1ff0ef;
		mem['h185] = 32'h00448793;
		mem['h186] = 32'h00f52023;
		mem['h187] = 32'h00a92223;
		mem['h188] = 32'h00400513;
		mem['h189] = 32'hc8dff0ef;
		mem['h18a] = 32'h00848793;
		mem['h18b] = 32'h00f52023;
		mem['h18c] = 32'h00a92423;
		mem['h18d] = 32'h00400513;
		mem['h18e] = 32'hc79ff0ef;
		mem['h18f] = 32'h00c48793;
		mem['h190] = 32'h00f52023;
		mem['h191] = 32'h00a92623;
		mem['h192] = 32'h00400513;
		mem['h193] = 32'hc65ff0ef;
		mem['h194] = 32'h01048793;
		mem['h195] = 32'h00f52023;
		mem['h196] = 32'h00a92823;
		mem['h197] = 32'h00400513;
		mem['h198] = 32'hc51ff0ef;
		mem['h199] = 32'h01448793;
		mem['h19a] = 32'h00f52023;
		mem['h19b] = 32'h00a92a23;
		mem['h19c] = 32'h00400513;
		mem['h19d] = 32'hc3dff0ef;
		mem['h19e] = 32'h01848793;
		mem['h19f] = 32'h00f52023;
		mem['h1a0] = 32'h00a92c23;
		mem['h1a1] = 32'h0129a023;
		mem['h1a2] = 32'h01c00513;
		mem['h1a3] = 32'hc25ff0ef;
		mem['h1a4] = 32'h00050913;
		mem['h1a5] = 32'h00400513;
		mem['h1a6] = 32'hc19ff0ef;
		mem['h1a7] = 32'h01c48793;
		mem['h1a8] = 32'h00f52023;
		mem['h1a9] = 32'h00a92023;
		mem['h1aa] = 32'h00400513;
		mem['h1ab] = 32'hc05ff0ef;
		mem['h1ac] = 32'h02048793;
		mem['h1ad] = 32'h00f52023;
		mem['h1ae] = 32'h00a92223;
		mem['h1af] = 32'h00400513;
		mem['h1b0] = 32'hbf1ff0ef;
		mem['h1b1] = 32'h02448793;
		mem['h1b2] = 32'h00f52023;
		mem['h1b3] = 32'h00a92423;
		mem['h1b4] = 32'h00400513;
		mem['h1b5] = 32'hbddff0ef;
		mem['h1b6] = 32'h02848793;
		mem['h1b7] = 32'h00f52023;
		mem['h1b8] = 32'h00a92623;
		mem['h1b9] = 32'h00400513;
		mem['h1ba] = 32'hbc9ff0ef;
		mem['h1bb] = 32'h02c48793;
		mem['h1bc] = 32'h00f52023;
		mem['h1bd] = 32'h00a92823;
		mem['h1be] = 32'h00400513;
		mem['h1bf] = 32'hbb5ff0ef;
		mem['h1c0] = 32'h03048793;
		mem['h1c1] = 32'h00f52023;
		mem['h1c2] = 32'h00a92a23;
		mem['h1c3] = 32'h00400513;
		mem['h1c4] = 32'hba1ff0ef;
		mem['h1c5] = 32'h03448793;
		mem['h1c6] = 32'h00f52023;
		mem['h1c7] = 32'h00a92c23;
		mem['h1c8] = 32'h0129a223;
		mem['h1c9] = 32'h01342023;
		mem['h1ca] = 32'h01000513;
		mem['h1cb] = 32'hb85ff0ef;
		mem['h1cc] = 32'h00050913;
		mem['h1cd] = 32'h00400513;
		mem['h1ce] = 32'hb79ff0ef;
		mem['h1cf] = 32'h03848793;
		mem['h1d0] = 32'h00f52023;
		mem['h1d1] = 32'h00a92023;
		mem['h1d2] = 32'h00400513;
		mem['h1d3] = 32'hb65ff0ef;
		mem['h1d4] = 32'h03c48793;
		mem['h1d5] = 32'h00f52023;
		mem['h1d6] = 32'h00a92223;
		mem['h1d7] = 32'h00400513;
		mem['h1d8] = 32'hb51ff0ef;
		mem['h1d9] = 32'h04048793;
		mem['h1da] = 32'h00f52023;
		mem['h1db] = 32'h00a92423;
		mem['h1dc] = 32'h00400513;
		mem['h1dd] = 32'hb3dff0ef;
		mem['h1de] = 32'h04448793;
		mem['h1df] = 32'h00f52023;
		mem['h1e0] = 32'h00a92623;
		mem['h1e1] = 32'h01242223;
		mem['h1e2] = 32'h00400513;
		mem['h1e3] = 32'hb25ff0ef;
		mem['h1e4] = 32'h04848793;
		mem['h1e5] = 32'h00f52023;
		mem['h1e6] = 32'h200009b7;
		mem['h1e7] = 32'h00a42423;
		mem['h1e8] = 32'h00c40a13;
		mem['h1e9] = 32'h04c48493;
		mem['h1ea] = 32'h07c98a93;
		mem['h1eb] = 32'h00c00513;
		mem['h1ec] = 32'hb01ff0ef;
		mem['h1ed] = 32'h00050913;
		mem['h1ee] = 32'h00400513;
		mem['h1ef] = 32'haf5ff0ef;
		mem['h1f0] = 32'h00952023;
		mem['h1f1] = 32'h00a92023;
		mem['h1f2] = 32'h00400513;
		mem['h1f3] = 32'hae5ff0ef;
		mem['h1f4] = 32'h00448793;
		mem['h1f5] = 32'h00f52023;
		mem['h1f6] = 32'h00a92223;
		mem['h1f7] = 32'h00400513;
		mem['h1f8] = 32'had1ff0ef;
		mem['h1f9] = 32'h00848793;
		mem['h1fa] = 32'h00f52023;
		mem['h1fb] = 32'h00a92423;
		mem['h1fc] = 32'h012a2023;
		mem['h1fd] = 32'h00c48493;
		mem['h1fe] = 32'h004a0a13;
		mem['h1ff] = 32'hfb5498e3;
		mem['h200] = 32'h00400513;
		mem['h201] = 32'haadff0ef;
		mem['h202] = 32'h00050913;
		mem['h203] = 32'h00400513;
		mem['h204] = 32'haa1ff0ef;
		mem['h205] = 32'h00952023;
		mem['h206] = 32'h00a92023;
		mem['h207] = 32'h01242e23;
		mem['h208] = 32'h00400513;
		mem['h209] = 32'ha8dff0ef;
		mem['h20a] = 32'h08098793;
		mem['h20b] = 32'h00f52023;
		mem['h20c] = 32'h02a42023;
		mem['h20d] = 32'h00400513;
		mem['h20e] = 32'ha79ff0ef;
		mem['h20f] = 32'h08498993;
		mem['h210] = 32'h01352023;
		mem['h211] = 32'h000014b7;
		mem['h212] = 32'h08c48593;
		mem['h213] = 32'h02a42223;
		mem['h214] = 32'h00040513;
		mem['h215] = 32'h91dff0ef;
		mem['h216] = 32'h000015b7;
		mem['h217] = 32'h0bc58593;
		mem['h218] = 32'h00040513;
		mem['h219] = 32'h90dff0ef;
		mem['h21a] = 32'h08c48593;
		mem['h21b] = 32'h00040513;
		mem['h21c] = 32'h901ff0ef;
		mem['h21d] = 32'h000015b7;
		mem['h21e] = 32'h0ec58593;
		mem['h21f] = 32'h00040513;
		mem['h220] = 32'h8f1ff0ef;
		mem['h221] = 32'h000015b7;
		mem['h222] = 32'h10458593;
		mem['h223] = 32'h00040513;
		mem['h224] = 32'h8e1ff0ef;
		mem['h225] = 32'h10000937;
		mem['h226] = 32'h00090593;
		mem['h227] = 32'h00040513;
		mem['h228] = 32'h915ff0ef;
		mem['h229] = 32'h000015b7;
		mem['h22a] = 32'h11c58593;
		mem['h22b] = 32'h00040513;
		mem['h22c] = 32'h00090493;
		mem['h22d] = 32'h8bdff0ef;
		mem['h22e] = 32'h00448593;
		mem['h22f] = 32'h00040513;
		mem['h230] = 32'h8f5ff0ef;
		mem['h231] = 32'h000015b7;
		mem['h232] = 32'h13858593;
		mem['h233] = 32'h00040513;
		mem['h234] = 32'h8a1ff0ef;
		mem['h235] = 32'h0084c583;
		mem['h236] = 32'h00040513;
		mem['h237] = 32'h100009b7;
		mem['h238] = 32'ha05ff0ef;
		mem['h239] = 32'h03a00593;
		mem['h23a] = 32'h00040513;
		mem['h23b] = 32'hf88ff0ef;
		mem['h23c] = 32'h0094c583;
		mem['h23d] = 32'h00040513;
		mem['h23e] = 32'h01898c93;
		mem['h23f] = 32'h9e9ff0ef;
		mem['h240] = 32'h03a00593;
		mem['h241] = 32'h00040513;
		mem['h242] = 32'hf6cff0ef;
		mem['h243] = 32'h00a4c583;
		mem['h244] = 32'h00040513;
		mem['h245] = 32'h00090a13;
		mem['h246] = 32'h9cdff0ef;
		mem['h247] = 32'h03a00593;
		mem['h248] = 32'h00040513;
		mem['h249] = 32'hf50ff0ef;
		mem['h24a] = 32'h00b4c583;
		mem['h24b] = 32'h00040513;
		mem['h24c] = 32'h01ec8a93;
		mem['h24d] = 32'h9b1ff0ef;
		mem['h24e] = 32'h03a00593;
		mem['h24f] = 32'h00040513;
		mem['h250] = 32'hf34ff0ef;
		mem['h251] = 32'h00c4c583;
		mem['h252] = 32'h00040513;
		mem['h253] = 32'h00ec8b13;
		mem['h254] = 32'h995ff0ef;
		mem['h255] = 32'h03a00593;
		mem['h256] = 32'h00040513;
		mem['h257] = 32'hf18ff0ef;
		mem['h258] = 32'h00d4c583;
		mem['h259] = 32'h00040513;
		mem['h25a] = 32'h97dff0ef;
		mem['h25b] = 32'h000015b7;
		mem['h25c] = 32'h15458593;
		mem['h25d] = 32'h00040513;
		mem['h25e] = 32'hff8ff0ef;
		mem['h25f] = 32'h00e48593;
		mem['h260] = 32'h00040513;
		mem['h261] = 32'h831ff0ef;
		mem['h262] = 32'h000015b7;
		mem['h263] = 32'h17058593;
		mem['h264] = 32'h00040513;
		mem['h265] = 32'hfdcff0ef;
		mem['h266] = 32'h0124c583;
		mem['h267] = 32'h00040513;
		mem['h268] = 32'h000014b7;
		mem['h269] = 32'hef8ff0ef;
		mem['h26a] = 32'h18c48593;
		mem['h26b] = 32'h00040513;
		mem['h26c] = 32'hfc0ff0ef;
		mem['h26d] = 32'h000015b7;
		mem['h26e] = 32'h19058593;
		mem['h26f] = 32'h00040513;
		mem['h270] = 32'hfb0ff0ef;
		mem['h271] = 32'h608c8793;
		mem['h272] = 32'h00f12423;
		mem['h273] = 32'h00f12623;
		mem['h274] = 32'h000c8023;
		mem['h275] = 32'h000c9123;
		mem['h276] = 32'h00042703;
		mem['h277] = 32'h00472703;
		mem['h278] = 32'h01872703;
		mem['h279] = 32'h00072703;
		mem['h27a] = 32'h00072703;
		mem['h27b] = 32'h00177713;
		mem['h27c] = 32'h10070c63;
		mem['h27d] = 32'h00042703;
		mem['h27e] = 32'h000c8b93;
		mem['h27f] = 32'h01898693;
		mem['h280] = 32'h00472703;
		mem['h281] = 32'h5f000513;
		mem['h282] = 32'h01072703;
		mem['h283] = 32'h00072703;
		mem['h284] = 32'h00072703;
		mem['h285] = 32'h00375713;
		mem['h286] = 32'h00777713;
		mem['h287] = 32'h00ec80a3;
		mem['h288] = 32'h00000713;
		mem['h289] = 32'h06e56263;
		mem['h28a] = 32'h00042603;
		mem['h28b] = 32'h00462603;
		mem['h28c] = 32'h00062603;
		mem['h28d] = 32'h00062603;
		mem['h28e] = 32'h00062603;
		mem['h28f] = 32'h00c6a423;
		mem['h290] = 32'h00042603;
		mem['h291] = 32'h00462603;
		mem['h292] = 32'h00462603;
		mem['h293] = 32'h00062603;
		mem['h294] = 32'h00062603;
		mem['h295] = 32'h00c6a623;
		mem['h296] = 32'h00042603;
		mem['h297] = 32'h00462603;
		mem['h298] = 32'h00862603;
		mem['h299] = 32'h00062603;
		mem['h29a] = 32'h00062603;
		mem['h29b] = 32'h00c6a823;
		mem['h29c] = 32'h00042603;
		mem['h29d] = 32'h00462603;
		mem['h29e] = 32'h00c62603;
		mem['h29f] = 32'h00062603;
		mem['h2a0] = 32'h00062603;
		mem['h2a1] = 32'h00c6aa23;
		mem['h2a2] = 32'h00042603;
		mem['h2a3] = 32'h01068693;
		mem['h2a4] = 32'h00462603;
		mem['h2a5] = 32'h01062603;
		mem['h2a6] = 32'h00062603;
		mem['h2a7] = 32'h00062603;
		mem['h2a8] = 32'h00f65613;
		mem['h2a9] = 32'h00167613;
		mem['h2aa] = 32'h06060c63;
		mem['h2ab] = 32'h00042683;
		mem['h2ac] = 32'h0046a683;
		mem['h2ad] = 32'h0106a683;
		mem['h2ae] = 32'h0006a683;
		mem['h2af] = 32'h0026d683;
		mem['h2b0] = 32'h0016f613;
		mem['h2b1] = 32'h00060863;
		mem['h2b2] = 32'h00170713;
		mem['h2b3] = 32'h0016d693;
		mem['h2b4] = 32'hff1ff06f;
		mem['h2b5] = 32'h60000693;
		mem['h2b6] = 32'h00e6f463;
		mem['h2b7] = 32'h60000713;
		mem['h2b8] = 32'h00eca223;
		mem['h2b9] = 32'h00042703;
		mem['h2ba] = 32'h00472703;
		mem['h2bb] = 32'h01472703;
		mem['h2bc] = 32'h00072683;
		mem['h2bd] = 32'h0006a703;
		mem['h2be] = 32'h00176713;
		mem['h2bf] = 32'h00e6a023;
		mem['h2c0] = 32'h004ca703;
		mem['h2c1] = 32'h04071063;
		mem['h2c2] = 32'h00842703;
		mem['h2c3] = 32'h00072683;
		mem['h2c4] = 32'h0006a703;
		mem['h2c5] = 32'hdff77713;
		mem['h2c6] = 32'h00e6a023;
		mem['h2c7] = 32'h3500006f;
		mem['h2c8] = 32'h00042603;
		mem['h2c9] = 32'h01070713;
		mem['h2ca] = 32'h00462603;
		mem['h2cb] = 32'h01462603;
		mem['h2cc] = 32'h00062583;
		mem['h2cd] = 32'h0005a603;
		mem['h2ce] = 32'h00166613;
		mem['h2cf] = 32'h00c5a023;
		mem['h2d0] = 32'hee5ff06f;
		mem['h2d1] = 32'h00842703;
		mem['h2d2] = 32'h00072683;
		mem['h2d3] = 32'h0006a703;
		mem['h2d4] = 32'h20076713;
		mem['h2d5] = 32'h00e6a023;
		mem['h2d6] = 32'h014ccc03;
		mem['h2d7] = 32'h00800713;
		mem['h2d8] = 32'h2eec1463;
		mem['h2d9] = 32'h015cc703;
		mem['h2da] = 32'h00600693;
		mem['h2db] = 32'h18d70663;
		mem['h2dc] = 32'h2c071c63;
		mem['h2dd] = 32'h016cc703;
		mem['h2de] = 32'h04000693;
		mem['h2df] = 32'h0f077713;
		mem['h2e0] = 32'h2cd71463;
		mem['h2e1] = 32'h01fcc683;
		mem['h2e2] = 32'h00100713;
		mem['h2e3] = 32'h2ae69e63;
		mem['h2e4] = 32'h000015b7;
		mem['h2e5] = 32'h1c058593;
		mem['h2e6] = 32'h00040513;
		mem['h2e7] = 32'hdd4ff0ef;
		mem['h2e8] = 32'h004cd583;
		mem['h2e9] = 32'h00040513;
		mem['h2ea] = 32'hcf4ff0ef;
		mem['h2eb] = 32'h18c48593;
		mem['h2ec] = 32'h00040513;
		mem['h2ed] = 32'hdbcff0ef;
		mem['h2ee] = 32'h00000713;
		mem['h2ef] = 32'h00400613;
		mem['h2f0] = 32'h00ea06b3;
		mem['h2f1] = 32'h026bc583;
		mem['h2f2] = 32'h0006c683;
		mem['h2f3] = 32'h26d59e63;
		mem['h2f4] = 32'h00170713;
		mem['h2f5] = 32'h001b8b93;
		mem['h2f6] = 32'hfec714e3;
		mem['h2f7] = 32'h02acc683;
		mem['h2f8] = 32'h00800713;
		mem['h2f9] = 32'h26e69263;
		mem['h2fa] = 32'h02bcc703;
		mem['h2fb] = 32'h24071e63;
		mem['h2fc] = 32'h001cc703;
		mem['h2fd] = 32'h00600613;
		mem['h2fe] = 32'h000b0593;
		mem['h2ff] = 32'h60ec8423;
		mem['h300] = 32'h00100713;
		mem['h301] = 32'h60ec85a3;
		mem['h302] = 32'h004ca703;
		mem['h303] = 32'h610c8513;
		mem['h304] = 32'h60eca623;
		mem['h305] = 32'h965ff0ef;
		mem['h306] = 32'h00600613;
		mem['h307] = 32'h008a0593;
		mem['h308] = 32'h616c8513;
		mem['h309] = 32'h955ff0ef;
		mem['h30a] = 32'h00450737;
		mem['h30b] = 32'h00870713;
		mem['h30c] = 32'h60ecae23;
		mem['h30d] = 32'h018cd703;
		mem['h30e] = 32'h00400613;
		mem['h30f] = 32'h00090593;
		mem['h310] = 32'h62ec9023;
		mem['h311] = 32'h62ac8513;
		mem['h312] = 32'h01ff0737;
		mem['h313] = 32'h62eca223;
		mem['h314] = 32'h620c9123;
		mem['h315] = 32'h620c9423;
		mem['h316] = 32'h921ff0ef;
		mem['h317] = 32'h00400613;
		mem['h318] = 32'h022c8593;
		mem['h319] = 32'h62ec8513;
		mem['h31a] = 32'h911ff0ef;
		mem['h31b] = 32'h01400593;
		mem['h31c] = 32'h61ec8513;
		mem['h31d] = 32'hdb8ff0ef;
		mem['h31e] = 32'h00851713;
		mem['h31f] = 32'h00855513;
		mem['h320] = 32'h00a76533;
		mem['h321] = 32'h02ecd703;
		mem['h322] = 32'h004ca603;
		mem['h323] = 32'h62ac9423;
		mem['h324] = 32'h62ec9b23;
		mem['h325] = 32'h030cd703;
		mem['h326] = 32'hfd660613;
		mem['h327] = 32'h032c8593;
		mem['h328] = 32'h63ac8513;
		mem['h329] = 32'h62ec9c23;
		mem['h32a] = 32'h620c9923;
		mem['h32b] = 32'h620c9a23;
		mem['h32c] = 32'h8c9ff0ef;
		mem['h32d] = 32'h004ca583;
		mem['h32e] = 32'h624b0513;
		mem['h32f] = 32'hfde58593;
		mem['h330] = 32'hd6cff0ef;
		mem['h331] = 32'h00851713;
		mem['h332] = 32'h00c12583;
		mem['h333] = 32'h00855513;
		mem['h334] = 32'h00a76533;
		mem['h335] = 32'h62ac9a23;
		mem['h336] = 32'h00040513;
		mem['h337] = 32'he64ff0ef;
		mem['h338] = 32'h000015b7;
		mem['h339] = 32'h1fc58593;
		mem['h33a] = 32'h00040513;
		mem['h33b] = 32'hc84ff0ef;
		mem['h33c] = 32'h004cd583;
		mem['h33d] = 32'h1400006f;
		mem['h33e] = 32'h000017b7;
		mem['h33f] = 32'h1d478593;
		mem['h340] = 32'h00040513;
		mem['h341] = 32'hc6cff0ef;
		mem['h342] = 32'h004cd583;
		mem['h343] = 32'h00040513;
		mem['h344] = 32'hb8cff0ef;
		mem['h345] = 32'h18c48593;
		mem['h346] = 32'h00040513;
		mem['h347] = 32'hc54ff0ef;
		mem['h348] = 32'h017cc683;
		mem['h349] = 32'h00100713;
		mem['h34a] = 32'h12e69063;
		mem['h34b] = 32'h018cc703;
		mem['h34c] = 32'h11871c63;
		mem['h34d] = 32'h016cc703;
		mem['h34e] = 32'h019cc683;
		mem['h34f] = 32'h00d76733;
		mem['h350] = 32'h0ff77713;
		mem['h351] = 32'h10071263;
		mem['h352] = 32'h00400613;
		mem['h353] = 32'h00ea06b3;
		mem['h354] = 32'h02ebc583;
		mem['h355] = 32'h0006c683;
		mem['h356] = 32'h0ed59863;
		mem['h357] = 32'h00170713;
		mem['h358] = 32'h001b8b93;
		mem['h359] = 32'hfec714e3;
		mem['h35a] = 32'h01ccc703;
		mem['h35b] = 32'h001cc683;
		mem['h35c] = 32'h0c071c63;
		mem['h35d] = 32'h01dcc703;
		mem['h35e] = 32'h00100613;
		mem['h35f] = 32'h0cc71663;
		mem['h360] = 32'h60ec85a3;
		mem['h361] = 32'h00600613;
		mem['h362] = 32'h02a00713;
		mem['h363] = 32'h000a8593;
		mem['h364] = 32'h610c8513;
		mem['h365] = 32'h60dc8423;
		mem['h366] = 32'h60eca623;
		mem['h367] = 32'hfdcff0ef;
		mem['h368] = 32'h008a0593;
		mem['h369] = 32'h00600613;
		mem['h36a] = 32'h616c8513;
		mem['h36b] = 32'hfccff0ef;
		mem['h36c] = 32'h01000737;
		mem['h36d] = 32'h60870713;
		mem['h36e] = 32'h60ecae23;
		mem['h36f] = 32'h04060737;
		mem['h370] = 32'h100007b7;
		mem['h371] = 32'h00870713;
		mem['h372] = 32'h00878593;
		mem['h373] = 32'h62eca023;
		mem['h374] = 32'h00600613;
		mem['h375] = 32'h20000713;
		mem['h376] = 32'h626c8513;
		mem['h377] = 32'h62ec9223;
		mem['h378] = 32'hf98ff0ef;
		mem['h379] = 32'h00400613;
		mem['h37a] = 32'h00090593;
		mem['h37b] = 32'h62cc8513;
		mem['h37c] = 32'hf88ff0ef;
		mem['h37d] = 32'h00600613;
		mem['h37e] = 32'h000a8593;
		mem['h37f] = 32'h630c8513;
		mem['h380] = 32'hf78ff0ef;
		mem['h381] = 32'h00400613;
		mem['h382] = 32'h024c8593;
		mem['h383] = 32'h636c8513;
		mem['h384] = 32'hf68ff0ef;
		mem['h385] = 32'h00812583;
		mem['h386] = 32'h00040513;
		mem['h387] = 32'hd24ff0ef;
		mem['h388] = 32'h000017b7;
		mem['h389] = 32'h1e878593;
		mem['h38a] = 32'h00040513;
		mem['h38b] = 32'hb44ff0ef;
		mem['h38c] = 32'h60ccd583;
		mem['h38d] = 32'h00040513;
		mem['h38e] = 32'ha64ff0ef;
		mem['h38f] = 32'h18c48593;
		mem['h390] = 32'h00040513;
		mem['h391] = 32'hb2cff0ef;
		mem['h392] = 32'h001cc683;
		mem['h393] = 32'h00100713;
		mem['h394] = 32'h0ee69a63;
		mem['h395] = 32'h00200713;
		mem['h396] = 32'h00ec8023;
		mem['h397] = 32'h00dc81a3;
		mem['h398] = 32'h01898593;
		mem['h399] = 32'h00040513;
		mem['h39a] = 32'hcd8ff0ef;
		mem['h39b] = 32'h00442703;
		mem['h39c] = 32'h00072703;
		mem['h39d] = 32'h00072703;
		mem['h39e] = 32'h00072583;
		mem['h39f] = 32'hb405dae3;
		mem['h3a0] = 32'h0ff5f713;
		mem['h3a1] = 32'h01200693;
		mem['h3a2] = 32'hb4d704e3;
		mem['h3a3] = 32'h01010b93;
		mem['h3a4] = 32'h00000c13;
		mem['h3a5] = 32'h00800d13;
		mem['h3a6] = 32'h07f00d93;
		mem['h3a7] = 32'h0ff5f593;
		mem['h3a8] = 32'h00bb8023;
		mem['h3a9] = 32'h00a00793;
		mem['h3aa] = 32'h02f58263;
		mem['h3ab] = 32'h00d00793;
		mem['h3ac] = 32'h0af59463;
		mem['h3ad] = 32'h00d00593;
		mem['h3ae] = 32'h00040513;
		mem['h3af] = 32'h9b8ff0ef;
		mem['h3b0] = 32'h00a00593;
		mem['h3b1] = 32'h00040513;
		mem['h3b2] = 32'h9acff0ef;
		mem['h3b3] = 32'h000b8023;
		mem['h3b4] = 32'h0ffc7c13;
		mem['h3b5] = 32'hae0c0ee3;
		mem['h3b6] = 32'h000015b7;
		mem['h3b7] = 32'h00040513;
		mem['h3b8] = 32'h21058593;
		mem['h3b9] = 32'ha8cff0ef;
		mem['h3ba] = 32'h01010593;
		mem['h3bb] = 32'h00040513;
		mem['h3bc] = 32'ha80ff0ef;
		mem['h3bd] = 32'h18c48593;
		mem['h3be] = 32'h00040513;
		mem['h3bf] = 32'ha74ff0ef;
		mem['h3c0] = 32'h000015b7;
		mem['h3c1] = 32'h00040513;
		mem['h3c2] = 32'h21c58593;
		mem['h3c3] = 32'ha64ff0ef;
		mem['h3c4] = 32'h000c0593;
		mem['h3c5] = 32'h00040513;
		mem['h3c6] = 32'h984ff0ef;
		mem['h3c7] = 32'h18c48593;
		mem['h3c8] = 32'h00040513;
		mem['h3c9] = 32'ha4cff0ef;
		mem['h3ca] = 32'h01014583;
		mem['h3cb] = 32'h00040513;
		mem['h3cc] = 32'hbb4ff0ef;
		mem['h3cd] = 32'h18c48593;
		mem['h3ce] = 32'h00040513;
		mem['h3cf] = 32'ha34ff0ef;
		mem['h3d0] = 32'ha91ff06f;
		mem['h3d1] = 32'h00200613;
		mem['h3d2] = 32'hf2c692e3;
		mem['h3d3] = 32'h00ec8023;
		mem['h3d4] = 32'h00ec81a3;
		mem['h3d5] = 32'hf0dff06f;
		mem['h3d6] = 32'h01a58463;
		mem['h3d7] = 32'h05b59a63;
		mem['h3d8] = 32'h020c0863;
		mem['h3d9] = 32'h00800593;
		mem['h3da] = 32'h00040513;
		mem['h3db] = 32'h908ff0ef;
		mem['h3dc] = 32'h02000593;
		mem['h3dd] = 32'h00040513;
		mem['h3de] = 32'h8fcff0ef;
		mem['h3df] = 32'h00800593;
		mem['h3e0] = 32'h00040513;
		mem['h3e1] = 32'hfffb8b93;
		mem['h3e2] = 32'hfffc0c13;
		mem['h3e3] = 32'h8e8ff0ef;
		mem['h3e4] = 32'h00442603;
		mem['h3e5] = 32'h00062603;
		mem['h3e6] = 32'h00062603;
		mem['h3e7] = 32'h00062583;
		mem['h3e8] = 32'hfe05d8e3;
		mem['h3e9] = 32'h01f00793;
		mem['h3ea] = 32'heefc1ae3;
		mem['h3eb] = 32'hf21ff06f;
		mem['h3ec] = 32'h00040513;
		mem['h3ed] = 32'h8c0ff0ef;
		mem['h3ee] = 32'h001b8b93;
		mem['h3ef] = 32'h001c0c13;
		mem['h3f0] = 32'hfd1ff06f;
		mem['h3f1] = 32'h06054063;
		mem['h3f2] = 32'h0605c663;
		mem['h3f3] = 32'h00058613;
		mem['h3f4] = 32'h00050593;
		mem['h3f5] = 32'hfff00513;
		mem['h3f6] = 32'h02060c63;
		mem['h3f7] = 32'h00100693;
		mem['h3f8] = 32'h00b67a63;
		mem['h3f9] = 32'h00c05863;
		mem['h3fa] = 32'h00161613;
		mem['h3fb] = 32'h00169693;
		mem['h3fc] = 32'hfeb66ae3;
		mem['h3fd] = 32'h00000513;
		mem['h3fe] = 32'h00c5e663;
		mem['h3ff] = 32'h40c585b3;
		mem['h400] = 32'h00d56533;
		mem['h401] = 32'h0016d693;
		mem['h402] = 32'h00165613;
		mem['h403] = 32'hfe0696e3;
		mem['h404] = 32'h00008067;
		mem['h405] = 32'h00008293;
		mem['h406] = 32'hfb5ff0ef;
		mem['h407] = 32'h00058513;
		mem['h408] = 32'h00028067;
		mem['h409] = 32'h40a00533;
		mem['h40a] = 32'h0005d863;
		mem['h40b] = 32'h40b005b3;
		mem['h40c] = 32'hf9dff06f;
		mem['h40d] = 32'h40b005b3;
		mem['h40e] = 32'h00008293;
		mem['h40f] = 32'hf91ff0ef;
		mem['h410] = 32'h40a00533;
		mem['h411] = 32'h00028067;
		mem['h412] = 32'h00008293;
		mem['h413] = 32'h0005ca63;
		mem['h414] = 32'h00054c63;
		mem['h415] = 32'hf79ff0ef;
		mem['h416] = 32'h00058513;
		mem['h417] = 32'h00028067;
		mem['h418] = 32'h40b005b3;
		mem['h419] = 32'hfe0558e3;
		mem['h41a] = 32'h40a00533;
		mem['h41b] = 32'hf61ff0ef;
		mem['h41c] = 32'h40b00533;
		mem['h41d] = 32'h00028067;
		mem['h41e] = 32'h33323130;
		mem['h41f] = 32'h37363534;
		mem['h420] = 32'h42413938;
		mem['h421] = 32'h46454443;
		mem['h422] = 32'h00000000;
		mem['h423] = 32'h3d3d3d3d;
		mem['h424] = 32'h3d3d3d3d;
		mem['h425] = 32'h3d3d3d3d;
		mem['h426] = 32'h3d3d3d3d;
		mem['h427] = 32'h3d3d3d3d;
		mem['h428] = 32'h3d3d3d3d;
		mem['h429] = 32'h3d3d3d3d;
		mem['h42a] = 32'h3d3d3d3d;
		mem['h42b] = 32'h3d3d3d3d;
		mem['h42c] = 32'h3d3d3d3d;
		mem['h42d] = 32'h0a0d3d3d;
		mem['h42e] = 32'h00000000;
		mem['h42f] = 32'h20202020;
		mem['h430] = 32'h57202020;
		mem['h431] = 32'h47657269;
		mem['h432] = 32'h64726175;
		mem['h433] = 32'h47504620;
		mem['h434] = 32'h79622041;
		mem['h435] = 32'h69684320;
		mem['h436] = 32'h6843696c;
		mem['h437] = 32'h20737069;
		mem['h438] = 32'h20202020;
		mem['h439] = 32'h0a0d2020;
		mem['h43a] = 32'h00000000;
		mem['h43b] = 32'h7774654e;
		mem['h43c] = 32'h206b726f;
		mem['h43d] = 32'h666e6f63;
		mem['h43e] = 32'h72756769;
		mem['h43f] = 32'h6f697461;
		mem['h440] = 32'h000a0d6e;
		mem['h441] = 32'h49202d2d;
		mem['h442] = 32'h64612050;
		mem['h443] = 32'h73657264;
		mem['h444] = 32'h20203a73;
		mem['h445] = 32'h20202020;
		mem['h446] = 32'h00002020;
		mem['h447] = 32'h2d2d0a0d;
		mem['h448] = 32'h62755320;
		mem['h449] = 32'h2074656e;
		mem['h44a] = 32'h6b73616d;
		mem['h44b] = 32'h2020203a;
		mem['h44c] = 32'h20202020;
		mem['h44d] = 32'h00000000;
		mem['h44e] = 32'h2d2d0a0d;
		mem['h44f] = 32'h43414d20;
		mem['h450] = 32'h64646120;
		mem['h451] = 32'h73736572;
		mem['h452] = 32'h2020203a;
		mem['h453] = 32'h20202020;
		mem['h454] = 32'h00000000;
		mem['h455] = 32'h2d2d0a0d;
		mem['h456] = 32'h66654420;
		mem['h457] = 32'h746c7561;
		mem['h458] = 32'h74616720;
		mem['h459] = 32'h79617765;
		mem['h45a] = 32'h2020203a;
		mem['h45b] = 32'h00000000;
		mem['h45c] = 32'h2d2d0a0d;
		mem['h45d] = 32'h66654420;
		mem['h45e] = 32'h746c7561;
		mem['h45f] = 32'h746e6920;
		mem['h460] = 32'h61667265;
		mem['h461] = 32'h203a6563;
		mem['h462] = 32'h00000000;
		mem['h463] = 32'h00000a0d;
		mem['h464] = 32'h2d2d2d2d;
		mem['h465] = 32'h2d2d2d2d;
		mem['h466] = 32'h2d2d2d2d;
		mem['h467] = 32'h2d2d2d2d;
		mem['h468] = 32'h2d2d2d2d;
		mem['h469] = 32'h2d2d2d2d;
		mem['h46a] = 32'h2d2d2d2d;
		mem['h46b] = 32'h2d2d2d2d;
		mem['h46c] = 32'h2d2d2d2d;
		mem['h46d] = 32'h2d2d2d2d;
		mem['h46e] = 32'h0a0d2d2d;
		mem['h46f] = 32'h00000000;
		mem['h470] = 32'h4e203c3c;
		mem['h471] = 32'h505f5445;
		mem['h472] = 32'h4f544f52;
		mem['h473] = 32'h4d43495f;
		mem['h474] = 32'h00203a50;
		mem['h475] = 32'h4e203c3c;
		mem['h476] = 32'h505f5445;
		mem['h477] = 32'h4f544f52;
		mem['h478] = 32'h5052415f;
		mem['h479] = 32'h0000203a;
		mem['h47a] = 32'h4e203e3e;
		mem['h47b] = 32'h505f5445;
		mem['h47c] = 32'h4f544f52;
		mem['h47d] = 32'h5052415f;
		mem['h47e] = 32'h0000203a;
		mem['h47f] = 32'h4e203e3e;
		mem['h480] = 32'h505f5445;
		mem['h481] = 32'h4f544f52;
		mem['h482] = 32'h4d43495f;
		mem['h483] = 32'h00203a50;
		mem['h484] = 32'h65636552;
		mem['h485] = 32'h64657669;
		mem['h486] = 32'h0000203a;
		mem['h487] = 32'h65636552;
		mem['h488] = 32'h64657669;
		mem['h489] = 32'h6e656c20;
		mem['h48a] = 32'h3a687467;
		mem['h48b] = 32'h00000020;
		mem['h48c] = 32'h6301a8c0;
		mem['h48d] = 32'h00ffffff;
		mem['h48e] = 32'haecccaca;
		mem['h48f] = 32'ha8c00100;
		mem['h490] = 32'h0001fe01;
		mem['h491] = 32'h00000000;
	end
	always @(posedge clk) begin
		rdat <= mem[raddr_int];
		if (we == 1'b1)
			mem[waddr_int] <= wdat;
	end
	always @(negedge arst_n or posedge clk)
		if (arst_n == 1'b0)
			rrdy <= 1'sb0;
		else
			rrdy <= rvld & ~rrdy;
endmodule