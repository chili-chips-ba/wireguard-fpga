-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.8297583002692854]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 2
entity VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_1CLK_5470451a is
port(
 clk : in std_logic;
 ref_toks_0 : in chacha20_state;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out unsigned(31 downto 0));
end VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_1CLK_5470451a;
architecture arch of VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_1CLK_5470451a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 1;
-- All of the wires/regs in function
-- Stage 0
-- Each function instance gets signals
-- uint32_mux16[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9]
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel : unsigned(3 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15 : unsigned(31 downto 0);
signal uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output : unsigned(31 downto 0);

function uint4_uint4_0( inp : unsigned;
 x : unsigned) return unsigned is

  --variable inp : unsigned(3 downto 0);
  --variable x : unsigned(3 downto 0);
  variable intermediate : unsigned(3 downto 0);
  variable return_output : unsigned(3 downto 0);

begin

    intermediate := (others => '0');
    intermediate(3 downto 0) := unsigned(inp);
    intermediate(3 downto 0) := x;
    
    return_output := intermediate(3 downto 0) ;
    
    return return_output;

end function;


begin

-- SUBMODULE INSTANCES 
-- uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9 : 1 clocks latency
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9 : entity work.uint32_mux16_1CLK_093fbfab port map (
clk,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15,
uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 ref_toks_0,
 var_dim_0,
 -- Registers
 -- Stage 0
 -- All submodule outputs
 uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_ref_toks_0 : chacha20_state;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : unsigned(31 downto 0);
 variable VAR_base : chacha20_state;
 variable VAR_ref_0 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l16_c10_a0fe_return_output : unsigned(31 downto 0);
 variable VAR_ref_1 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l18_c10_6d34_return_output : unsigned(31 downto 0);
 variable VAR_ref_2 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l20_c10_88d2_return_output : unsigned(31 downto 0);
 variable VAR_ref_3 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l22_c10_772d_return_output : unsigned(31 downto 0);
 variable VAR_ref_4 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l24_c10_39f2_return_output : unsigned(31 downto 0);
 variable VAR_ref_5 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l26_c10_da31_return_output : unsigned(31 downto 0);
 variable VAR_ref_6 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l28_c10_3480_return_output : unsigned(31 downto 0);
 variable VAR_ref_7 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l30_c10_44f7_return_output : unsigned(31 downto 0);
 variable VAR_ref_8 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l32_c10_4e3a_return_output : unsigned(31 downto 0);
 variable VAR_ref_9 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l34_c10_e7a0_return_output : unsigned(31 downto 0);
 variable VAR_ref_10 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l36_c11_e055_return_output : unsigned(31 downto 0);
 variable VAR_ref_11 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l38_c11_ff64_return_output : unsigned(31 downto 0);
 variable VAR_ref_12 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l40_c11_f3dd_return_output : unsigned(31 downto 0);
 variable VAR_ref_13 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l42_c11_c621_return_output : unsigned(31 downto 0);
 variable VAR_ref_14 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l44_c11_69e4_return_output : unsigned(31 downto 0);
 variable VAR_ref_15 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l46_c11_ac30_return_output : unsigned(31 downto 0);
 variable VAR_sel : unsigned(3 downto 0);
 variable VAR_uint4_uint4_0_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l50_c8_7b43_return_output : unsigned(3 downto 0);
 variable VAR_rv : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel : unsigned(3 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15 : unsigned(31 downto 0);
 variable VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output : unsigned(31 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     -- CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l18_c10_6d34] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l18_c10_6d34_return_output := VAR_ref_toks_0.state(1);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l28_c10_3480] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l28_c10_3480_return_output := VAR_ref_toks_0.state(6);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l32_c10_4e3a] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l32_c10_4e3a_return_output := VAR_ref_toks_0.state(8);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l34_c10_e7a0] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l34_c10_e7a0_return_output := VAR_ref_toks_0.state(9);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l22_c10_772d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l22_c10_772d_return_output := VAR_ref_toks_0.state(3);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l20_c10_88d2] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l20_c10_88d2_return_output := VAR_ref_toks_0.state(2);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l30_c10_44f7] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l30_c10_44f7_return_output := VAR_ref_toks_0.state(7);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l24_c10_39f2] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l24_c10_39f2_return_output := VAR_ref_toks_0.state(4);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l42_c11_c621] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l42_c11_c621_return_output := VAR_ref_toks_0.state(13);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l40_c11_f3dd] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l40_c11_f3dd_return_output := VAR_ref_toks_0.state(12);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l16_c10_a0fe] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l16_c10_a0fe_return_output := VAR_ref_toks_0.state(0);

     -- uint4_uint4_0[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l50_c8_7b43] LATENCY=0
     VAR_uint4_uint4_0_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l50_c8_7b43_return_output := uint4_uint4_0(
     to_unsigned(0, 4),
     VAR_var_dim_0);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l26_c10_da31] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l26_c10_da31_return_output := VAR_ref_toks_0.state(5);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l44_c11_69e4] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l44_c11_69e4_return_output := VAR_ref_toks_0.state(14);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l46_c11_ac30] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l46_c11_ac30_return_output := VAR_ref_toks_0.state(15);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l36_c11_e055] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l36_c11_e055_return_output := VAR_ref_toks_0.state(10);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l38_c11_ff64] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l38_c11_ff64_return_output := VAR_ref_toks_0.state(11);

     -- Submodule level 1
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l16_c10_a0fe_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l36_c11_e055_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l38_c11_ff64_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l40_c11_f3dd_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l42_c11_c621_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l44_c11_69e4_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l46_c11_ac30_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l18_c10_6d34_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l20_c10_88d2_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l22_c10_772d_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l24_c10_39f2_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l26_c10_da31_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l28_c10_3480_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l30_c10_44f7_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l32_c10_4e3a_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9 := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l34_c10_e7a0_return_output;
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel := VAR_uint4_uint4_0_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l50_c8_7b43_return_output;
     -- uint32_mux16[VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9] LATENCY=1
     -- Inputs
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_sel;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in0;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in1;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in2;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in3;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in4;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in5;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in6;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in7;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in8;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in9;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in10;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in11;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in12;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in13;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in14;
     uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15 <= VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_in15;

     -- Write to comb signals
   elsif STAGE = 1 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output := uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output;

     -- Submodule level 0
     VAR_return_output := VAR_uint32_mux16_VAR_REF_RD_uint32_t_chacha20_state_state_VAR_d41d_c_l53_c7_c3d9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
 end if;
end process;

end arch;
