-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 11
entity bytes_to_u320_t_0CLK_4bbc8984 is
port(
 bytes : in uint8_t_40;
 return_output : out u320_t);
end bytes_to_u320_t_0CLK_4bbc8984;
architecture arch of bytes_to_u320_t_0CLK_4bbc8984 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997]
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997]
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997]
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997]
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997]
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
signal FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);

function CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return uint8_t_array_8_t is
 
  variable base : uint8_t_array_8_t; 
  variable return_output : uint8_t_array_8_t;
begin
      base.data(0) := ref_toks_0;
      base.data(1) := ref_toks_1;
      base.data(2) := ref_toks_2;
      base.data(3) := ref_toks_3;
      base.data(4) := ref_toks_4;
      base.data(5) := ref_toks_5;
      base.data(6) := ref_toks_6;
      base.data(7) := ref_toks_7;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : 0 clocks latency
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : entity work.bytes_to_uint64_t_0CLK_36723c85 port map (
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes,
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : 0 clocks latency
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : entity work.bytes_to_uint64_t_0CLK_36723c85 port map (
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes,
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : 0 clocks latency
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : entity work.bytes_to_uint64_t_0CLK_36723c85 port map (
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes,
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : 0 clocks latency
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : entity work.bytes_to_uint64_t_0CLK_36723c85 port map (
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes,
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);

-- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : 0 clocks latency
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997 : entity work.bytes_to_uint64_t_0CLK_36723c85 port map (
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes,
FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 bytes,
 -- All submodule outputs
 FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
 FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
 FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
 FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
 FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_bytes : uint8_t_40;
 variable VAR_rv : u320_t;
 variable VAR_pos : unsigned(6 downto 0);
 variable VAR_field_pos : unsigned(6 downto 0);
 variable VAR_limbs_dim_0 : unsigned(2 downto 0);
 variable VAR_limbs_elem_bytes : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_0_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_1_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_2_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_3_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_4_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_5_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_6_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_7_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_8_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_9_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_10_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_11_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_12_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_13_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_14_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_15_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_16_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_17_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_18_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_19_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_20_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_21_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_22_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_23_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_24_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_25_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_26_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_27_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_28_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_29_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_30_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_31_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_32_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_33_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_34_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_35_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_36_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_37_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_38_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_39_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes : uint8_t_8;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_u320_t_bytes_t_h_l54_c12_966b_return_output : u320_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_bytes := bytes;

     -- Submodule level 0
     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_24_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_24_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(24);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_26_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_26_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(26);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_34_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_34_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(34);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_28_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_28_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(28);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_39_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_39_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(39);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_33_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_33_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(33);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_9_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_9_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(9);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_35_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_35_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(35);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_6_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_6_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(6);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_14_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_14_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(14);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_10_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_10_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(10);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_2_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_2_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(2);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_4_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_4_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(4);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_7_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_7_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(7);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_38_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_38_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(38);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_12_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_12_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(12);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_19_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_19_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(19);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_20_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_20_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(20);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_23_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_23_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(23);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_27_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_27_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(27);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_16_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_16_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(16);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_15_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_15_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(15);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_3_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_3_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(3);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_25_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_25_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(25);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_8_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_8_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(8);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_32_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_32_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(32);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_17_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_17_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(17);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_13_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_13_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(13);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_22_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_22_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(22);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_36_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_36_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(36);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_30_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_30_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(30);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_37_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_37_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(37);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_18_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_18_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(18);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_1_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_1_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(1);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_5_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_5_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(5);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_31_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_31_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(31);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_29_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_29_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(29);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_11_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_11_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(11);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_0_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_0_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(0);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_21_d41d[u320_t_bytes_t_h_l48_c40_1d0a] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_21_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output := VAR_bytes(21);

     -- Submodule level 1
     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58[u320_t_bytes_t_h_l51_c44_62ad] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_0_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_1_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_2_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_3_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_4_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_5_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_6_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_7_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58[u320_t_bytes_t_h_l51_c44_62ad] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_8_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_9_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_10_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_11_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_12_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_13_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_14_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_15_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58[u320_t_bytes_t_h_l51_c44_62ad] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_32_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_33_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_34_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_35_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_36_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_37_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_38_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_39_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58[u320_t_bytes_t_h_l51_c44_62ad] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_24_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_25_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_26_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_27_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_28_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_29_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_30_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_31_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output);

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58[u320_t_bytes_t_h_l51_c44_62ad] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output := CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_0_CONST_REF_RD_uint8_t_uint8_t_40_16_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_1_CONST_REF_RD_uint8_t_uint8_t_40_17_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_2_CONST_REF_RD_uint8_t_uint8_t_40_18_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_3_CONST_REF_RD_uint8_t_uint8_t_40_19_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_4_CONST_REF_RD_uint8_t_uint8_t_40_20_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_5_CONST_REF_RD_uint8_t_uint8_t_40_21_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_6_CONST_REF_RD_uint8_t_uint8_t_40_22_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_FOR_u320_t_bytes_t_h_l46_c2_5ec4_ITER_7_CONST_REF_RD_uint8_t_uint8_t_40_23_d41d_u320_t_bytes_t_h_l48_c40_1d0a_return_output);

     -- Submodule level 2
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes := VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output.data;
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes := VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output.data;
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes := VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output.data;
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes := VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output.data;
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes := VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_CONST_REF_RD_uint8_t_array_8_t_uint8_t_array_8_t_dd58_u320_t_bytes_t_h_l51_c44_62ad_return_output.data;
     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes <= VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output := FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output;

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes <= VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output := FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output;

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes <= VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output := FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output;

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes <= VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output := FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output;

     -- FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t[u320_t_bytes_t_h_l51_c26_a997] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes <= VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_bytes;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output := FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output;

     -- Submodule level 3
     -- CONST_REF_RD_u320_t_u320_t_4216[u320_t_bytes_t_h_l54_c12_966b] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_u320_t_bytes_t_h_l54_c12_966b_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_0_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_1_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_2_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_3_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output,
     VAR_FOR_u320_t_bytes_t_h_l44_c1_e4c5_ITER_4_bytes_to_uint64_t_u320_t_bytes_t_h_l51_c26_a997_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_u320_t_bytes_t_h_l54_c12_966b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
