-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.20810055865921787, 0.5921787709497207, 0.9762569832402235]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_3CLK_087b5579 is
port(
 clk : in std_logic;
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_3CLK_087b5579;
architecture arch of uint320_mul_3CLK_087b5579 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 3;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
-- Stage 1
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
-- Stage 2
signal REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_e005]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_b61a]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_c337]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_6d5f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_6bf0]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_1e2f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_9a58]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_ce9b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_2247]
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_fe92]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_287e]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_d308]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_acdd]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_af5b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_ecee]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_efb1]
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_8db2]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_2aa9]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_e444]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_f304]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_9121]
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_0af7]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_ca04]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_40d3]
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41]
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d2a3]
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005 : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_9ca18c4f port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809 : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_eec62983 port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right,
FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd : entity work.BIN_OP_PLUS_uint64_t_uint1_t_1CLK_9324e8e6 port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0f464748 port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right,
FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_ec635a74 port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2 : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0320092f port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right,
FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right,
FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : 0 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output);

-- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3 : 1 clocks latency
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_8f2211ba port map (
clk,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right,
FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- Registers
 -- Stage 0
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 -- Stage 1
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left,
 -- Stage 2
 REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output,
 FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_2909_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_2909_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_2909_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_2909_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3588_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_2909_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_33d1_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_15b2_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3588_DUPLICATE_3414_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3588_DUPLICATE_6312_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_37a2_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5e9d_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse := to_unsigned(0, 1);
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_2909] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_2909_return_output := u320_t_NULL.limbs(4);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_2909] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_2909_return_output := u320_t_NULL.limbs(2);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_2909] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_2909_return_output := u320_t_NULL.limbs(1);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_2909] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_2909_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_2909] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_2909_return_output := u320_t_NULL.limbs(0);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_2909_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_2909_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_2909_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_2909_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_2909_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_3588]_DUPLICATE_6312 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3588_DUPLICATE_6312_return_output := VAR_b.limbs(3);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_3588] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3588_return_output := VAR_b.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_3588]_DUPLICATE_3414 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3588_DUPLICATE_3414_return_output := VAR_b.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_3588]_DUPLICATE_29d2 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_33d1]_DUPLICATE_8b1c LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output := VAR_a.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_33d1]_DUPLICATE_37a2 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_37a2_return_output := VAR_a.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_33d1]_DUPLICATE_5a5c LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output := VAR_a.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_3588]_DUPLICATE_efbc LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output := VAR_b.limbs(0);

     -- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_33d1] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_33d1_return_output := VAR_a.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_33d1]_DUPLICATE_5e9d LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5e9d_return_output := VAR_a.limbs(3);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5a5c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3588_DUPLICATE_efbc_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_8b1c_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3588_DUPLICATE_29d2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_37a2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_37a2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_37a2_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3588_DUPLICATE_3414_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3588_DUPLICATE_3414_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3588_DUPLICATE_3414_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5e9d_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_33d1_DUPLICATE_5e9d_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3588_DUPLICATE_6312_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3588_DUPLICATE_6312_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3588_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_33d1_return_output;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_product_poly1305_h_l127_c22_94f8_0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_product_poly1305_h_l127_c22_94f8_0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_e005] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;

     -- Write to comb signals
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e005_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l132_c21_b405_return_output;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_b61a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_b61a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_c337] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_fe92] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe92_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_6d5f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_6d5f_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_6bf0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_287e] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_287e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_d308] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d308_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_1e2f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1e2f_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_8db2] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_9a58] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_acdd] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_right;

     -- Write to comb signals
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left := REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_acdd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_8db2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_af5b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_af5b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_ce9b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_2247] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_2aa9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_2aa9_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_e444] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_ecee] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ecee_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_e444_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_efb1] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_efb1_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_8e3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_0af7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0af7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l131_c13_48c0;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_f304] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b809] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l132_c21_b405] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_f304_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b809_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l132_c21_b405_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_high_poly1305_h_l134_c13_6b46;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX[poly1305_h_l134_c22_dd3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_cond;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iftrue;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_9121] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_9121_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_MUX_poly1305_h_l134_c22_dd3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_ca04] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output;

     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_ca04_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_high_poly1305_h_l134_c13_6b46;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_40d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_40d3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_low_poly1305_h_l133_c13_1414;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_0b41] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left := VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l131_c13_48c0;
     -- FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d2a3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_left;
     FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_right;

     -- Write to comb signals
     COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output := FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 := resize(VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d2a3_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_15b2] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_15b2_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414,
     VAR_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_15b2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_c337_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_6bf0_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_9a58_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     -- Stage 1
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_ce9b_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_2247_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_8e3f_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_5c01_ITER_4_FOR_poly1305_h_l123_c9_0ea6_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_0b41_left;
     -- Stage 2
     REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_0_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_1_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_2_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
     REG_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_5c01_ITER_3_FOR_poly1305_h_l123_c9_0ea6_ITER_0_low_poly1305_h_l133_c13_1414;
 end if;
end process;

end arch;
