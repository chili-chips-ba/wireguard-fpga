-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 1
entity print_aad_0CLK_fa355561 is
port(
 CLOCK_ENABLE : in unsigned(0 downto 0);
 aad : in uint8_t_32;
 aad_len : in unsigned(31 downto 0));
end print_aad_0CLK_fa355561;
architecture arch of print_aad_0CLK_fa355561 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814[chacha20poly1305_decrypt_tb_c_l42_c5_5814]
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31 : unsigned(7 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32 : unsigned(7 downto 0);


begin

-- SUBMODULE INSTANCES 
-- printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814 : entity work.printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31,
printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Inputs
 aad,
 aad_len)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_aad : uint8_t_32;
 variable VAR_aad_len : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_0_d41d_chacha20poly1305_decrypt_tb_c_l53_c9_f784_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_1_d41d_chacha20poly1305_decrypt_tb_c_l53_c17_ad97_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_2_d41d_chacha20poly1305_decrypt_tb_c_l53_c25_2390_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_3_d41d_chacha20poly1305_decrypt_tb_c_l53_c33_c5b4_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_4_d41d_chacha20poly1305_decrypt_tb_c_l54_c9_2fa0_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_5_d41d_chacha20poly1305_decrypt_tb_c_l54_c17_ab39_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_6_d41d_chacha20poly1305_decrypt_tb_c_l54_c25_edba_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_7_d41d_chacha20poly1305_decrypt_tb_c_l54_c33_1286_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_8_d41d_chacha20poly1305_decrypt_tb_c_l55_c9_2fa1_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_9_d41d_chacha20poly1305_decrypt_tb_c_l55_c17_a88f_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_10_d41d_chacha20poly1305_decrypt_tb_c_l55_c25_e597_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_11_d41d_chacha20poly1305_decrypt_tb_c_l55_c34_3217_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_12_d41d_chacha20poly1305_decrypt_tb_c_l56_c9_9a70_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_13_d41d_chacha20poly1305_decrypt_tb_c_l56_c18_7a86_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_14_d41d_chacha20poly1305_decrypt_tb_c_l56_c27_1a6e_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_15_d41d_chacha20poly1305_decrypt_tb_c_l56_c36_153a_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_16_d41d_chacha20poly1305_decrypt_tb_c_l57_c9_97c2_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_17_d41d_chacha20poly1305_decrypt_tb_c_l57_c18_2754_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_18_d41d_chacha20poly1305_decrypt_tb_c_l57_c27_17e8_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_19_d41d_chacha20poly1305_decrypt_tb_c_l57_c36_a361_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_20_d41d_chacha20poly1305_decrypt_tb_c_l58_c9_2d02_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_21_d41d_chacha20poly1305_decrypt_tb_c_l58_c18_b4c6_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_22_d41d_chacha20poly1305_decrypt_tb_c_l58_c27_dcb8_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_23_d41d_chacha20poly1305_decrypt_tb_c_l58_c36_bf9d_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_24_d41d_chacha20poly1305_decrypt_tb_c_l59_c9_bf41_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_25_d41d_chacha20poly1305_decrypt_tb_c_l59_c18_e6ef_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_26_d41d_chacha20poly1305_decrypt_tb_c_l59_c27_04ee_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_27_d41d_chacha20poly1305_decrypt_tb_c_l59_c36_3e06_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_28_d41d_chacha20poly1305_decrypt_tb_c_l60_c9_6ad8_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_29_d41d_chacha20poly1305_decrypt_tb_c_l60_c18_76e3_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_30_d41d_chacha20poly1305_decrypt_tb_c_l60_c27_7fac_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31 : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_32_31_d41d_chacha20poly1305_decrypt_tb_c_l60_c36_5acc_return_output : unsigned(7 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32 : unsigned(7 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;
     -- Mux in inputs
     VAR_aad := aad;
     VAR_aad_len := aad_len;

     -- Submodule level 0
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0 := VAR_aad_len;
     -- CONST_REF_RD_uint8_t_uint8_t_32_5_d41d[chacha20poly1305_decrypt_tb_c_l54_c17_ab39] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_5_d41d_chacha20poly1305_decrypt_tb_c_l54_c17_ab39_return_output := VAR_aad(5);

     -- CONST_REF_RD_uint8_t_uint8_t_32_28_d41d[chacha20poly1305_decrypt_tb_c_l60_c9_6ad8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_28_d41d_chacha20poly1305_decrypt_tb_c_l60_c9_6ad8_return_output := VAR_aad(28);

     -- CONST_REF_RD_uint8_t_uint8_t_32_2_d41d[chacha20poly1305_decrypt_tb_c_l53_c25_2390] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_2_d41d_chacha20poly1305_decrypt_tb_c_l53_c25_2390_return_output := VAR_aad(2);

     -- CONST_REF_RD_uint8_t_uint8_t_32_4_d41d[chacha20poly1305_decrypt_tb_c_l54_c9_2fa0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_4_d41d_chacha20poly1305_decrypt_tb_c_l54_c9_2fa0_return_output := VAR_aad(4);

     -- CONST_REF_RD_uint8_t_uint8_t_32_29_d41d[chacha20poly1305_decrypt_tb_c_l60_c18_76e3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_29_d41d_chacha20poly1305_decrypt_tb_c_l60_c18_76e3_return_output := VAR_aad(29);

     -- CONST_REF_RD_uint8_t_uint8_t_32_1_d41d[chacha20poly1305_decrypt_tb_c_l53_c17_ad97] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_1_d41d_chacha20poly1305_decrypt_tb_c_l53_c17_ad97_return_output := VAR_aad(1);

     -- CONST_REF_RD_uint8_t_uint8_t_32_22_d41d[chacha20poly1305_decrypt_tb_c_l58_c27_dcb8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_22_d41d_chacha20poly1305_decrypt_tb_c_l58_c27_dcb8_return_output := VAR_aad(22);

     -- CONST_REF_RD_uint8_t_uint8_t_32_17_d41d[chacha20poly1305_decrypt_tb_c_l57_c18_2754] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_17_d41d_chacha20poly1305_decrypt_tb_c_l57_c18_2754_return_output := VAR_aad(17);

     -- CONST_REF_RD_uint8_t_uint8_t_32_16_d41d[chacha20poly1305_decrypt_tb_c_l57_c9_97c2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_16_d41d_chacha20poly1305_decrypt_tb_c_l57_c9_97c2_return_output := VAR_aad(16);

     -- CONST_REF_RD_uint8_t_uint8_t_32_18_d41d[chacha20poly1305_decrypt_tb_c_l57_c27_17e8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_18_d41d_chacha20poly1305_decrypt_tb_c_l57_c27_17e8_return_output := VAR_aad(18);

     -- CONST_REF_RD_uint8_t_uint8_t_32_8_d41d[chacha20poly1305_decrypt_tb_c_l55_c9_2fa1] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_8_d41d_chacha20poly1305_decrypt_tb_c_l55_c9_2fa1_return_output := VAR_aad(8);

     -- CONST_REF_RD_uint8_t_uint8_t_32_15_d41d[chacha20poly1305_decrypt_tb_c_l56_c36_153a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_15_d41d_chacha20poly1305_decrypt_tb_c_l56_c36_153a_return_output := VAR_aad(15);

     -- CONST_REF_RD_uint8_t_uint8_t_32_21_d41d[chacha20poly1305_decrypt_tb_c_l58_c18_b4c6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_21_d41d_chacha20poly1305_decrypt_tb_c_l58_c18_b4c6_return_output := VAR_aad(21);

     -- CONST_REF_RD_uint8_t_uint8_t_32_13_d41d[chacha20poly1305_decrypt_tb_c_l56_c18_7a86] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_13_d41d_chacha20poly1305_decrypt_tb_c_l56_c18_7a86_return_output := VAR_aad(13);

     -- CONST_REF_RD_uint8_t_uint8_t_32_12_d41d[chacha20poly1305_decrypt_tb_c_l56_c9_9a70] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_12_d41d_chacha20poly1305_decrypt_tb_c_l56_c9_9a70_return_output := VAR_aad(12);

     -- CONST_REF_RD_uint8_t_uint8_t_32_25_d41d[chacha20poly1305_decrypt_tb_c_l59_c18_e6ef] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_25_d41d_chacha20poly1305_decrypt_tb_c_l59_c18_e6ef_return_output := VAR_aad(25);

     -- CONST_REF_RD_uint8_t_uint8_t_32_6_d41d[chacha20poly1305_decrypt_tb_c_l54_c25_edba] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_6_d41d_chacha20poly1305_decrypt_tb_c_l54_c25_edba_return_output := VAR_aad(6);

     -- CONST_REF_RD_uint8_t_uint8_t_32_30_d41d[chacha20poly1305_decrypt_tb_c_l60_c27_7fac] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_30_d41d_chacha20poly1305_decrypt_tb_c_l60_c27_7fac_return_output := VAR_aad(30);

     -- CONST_REF_RD_uint8_t_uint8_t_32_27_d41d[chacha20poly1305_decrypt_tb_c_l59_c36_3e06] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_27_d41d_chacha20poly1305_decrypt_tb_c_l59_c36_3e06_return_output := VAR_aad(27);

     -- CONST_REF_RD_uint8_t_uint8_t_32_9_d41d[chacha20poly1305_decrypt_tb_c_l55_c17_a88f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_9_d41d_chacha20poly1305_decrypt_tb_c_l55_c17_a88f_return_output := VAR_aad(9);

     -- CONST_REF_RD_uint8_t_uint8_t_32_23_d41d[chacha20poly1305_decrypt_tb_c_l58_c36_bf9d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_23_d41d_chacha20poly1305_decrypt_tb_c_l58_c36_bf9d_return_output := VAR_aad(23);

     -- CONST_REF_RD_uint8_t_uint8_t_32_31_d41d[chacha20poly1305_decrypt_tb_c_l60_c36_5acc] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_31_d41d_chacha20poly1305_decrypt_tb_c_l60_c36_5acc_return_output := VAR_aad(31);

     -- CONST_REF_RD_uint8_t_uint8_t_32_3_d41d[chacha20poly1305_decrypt_tb_c_l53_c33_c5b4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_3_d41d_chacha20poly1305_decrypt_tb_c_l53_c33_c5b4_return_output := VAR_aad(3);

     -- CONST_REF_RD_uint8_t_uint8_t_32_24_d41d[chacha20poly1305_decrypt_tb_c_l59_c9_bf41] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_24_d41d_chacha20poly1305_decrypt_tb_c_l59_c9_bf41_return_output := VAR_aad(24);

     -- CONST_REF_RD_uint8_t_uint8_t_32_14_d41d[chacha20poly1305_decrypt_tb_c_l56_c27_1a6e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_14_d41d_chacha20poly1305_decrypt_tb_c_l56_c27_1a6e_return_output := VAR_aad(14);

     -- CONST_REF_RD_uint8_t_uint8_t_32_7_d41d[chacha20poly1305_decrypt_tb_c_l54_c33_1286] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_7_d41d_chacha20poly1305_decrypt_tb_c_l54_c33_1286_return_output := VAR_aad(7);

     -- CONST_REF_RD_uint8_t_uint8_t_32_20_d41d[chacha20poly1305_decrypt_tb_c_l58_c9_2d02] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_20_d41d_chacha20poly1305_decrypt_tb_c_l58_c9_2d02_return_output := VAR_aad(20);

     -- CONST_REF_RD_uint8_t_uint8_t_32_26_d41d[chacha20poly1305_decrypt_tb_c_l59_c27_04ee] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_26_d41d_chacha20poly1305_decrypt_tb_c_l59_c27_04ee_return_output := VAR_aad(26);

     -- CONST_REF_RD_uint8_t_uint8_t_32_0_d41d[chacha20poly1305_decrypt_tb_c_l53_c9_f784] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_0_d41d_chacha20poly1305_decrypt_tb_c_l53_c9_f784_return_output := VAR_aad(0);

     -- CONST_REF_RD_uint8_t_uint8_t_32_11_d41d[chacha20poly1305_decrypt_tb_c_l55_c34_3217] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_11_d41d_chacha20poly1305_decrypt_tb_c_l55_c34_3217_return_output := VAR_aad(11);

     -- CONST_REF_RD_uint8_t_uint8_t_32_10_d41d[chacha20poly1305_decrypt_tb_c_l55_c25_e597] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_10_d41d_chacha20poly1305_decrypt_tb_c_l55_c25_e597_return_output := VAR_aad(10);

     -- CONST_REF_RD_uint8_t_uint8_t_32_19_d41d[chacha20poly1305_decrypt_tb_c_l57_c36_a361] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_32_19_d41d_chacha20poly1305_decrypt_tb_c_l57_c36_a361_return_output := VAR_aad(19);

     -- Submodule level 1
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_0_d41d_chacha20poly1305_decrypt_tb_c_l53_c9_f784_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_10_d41d_chacha20poly1305_decrypt_tb_c_l55_c25_e597_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_11_d41d_chacha20poly1305_decrypt_tb_c_l55_c34_3217_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_12_d41d_chacha20poly1305_decrypt_tb_c_l56_c9_9a70_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_13_d41d_chacha20poly1305_decrypt_tb_c_l56_c18_7a86_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_14_d41d_chacha20poly1305_decrypt_tb_c_l56_c27_1a6e_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_15_d41d_chacha20poly1305_decrypt_tb_c_l56_c36_153a_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_16_d41d_chacha20poly1305_decrypt_tb_c_l57_c9_97c2_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_17_d41d_chacha20poly1305_decrypt_tb_c_l57_c18_2754_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_18_d41d_chacha20poly1305_decrypt_tb_c_l57_c27_17e8_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_19_d41d_chacha20poly1305_decrypt_tb_c_l57_c36_a361_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_1_d41d_chacha20poly1305_decrypt_tb_c_l53_c17_ad97_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_20_d41d_chacha20poly1305_decrypt_tb_c_l58_c9_2d02_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_21_d41d_chacha20poly1305_decrypt_tb_c_l58_c18_b4c6_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_22_d41d_chacha20poly1305_decrypt_tb_c_l58_c27_dcb8_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_23_d41d_chacha20poly1305_decrypt_tb_c_l58_c36_bf9d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_24_d41d_chacha20poly1305_decrypt_tb_c_l59_c9_bf41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_25_d41d_chacha20poly1305_decrypt_tb_c_l59_c18_e6ef_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_26_d41d_chacha20poly1305_decrypt_tb_c_l59_c27_04ee_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_27_d41d_chacha20poly1305_decrypt_tb_c_l59_c36_3e06_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_28_d41d_chacha20poly1305_decrypt_tb_c_l60_c9_6ad8_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_29_d41d_chacha20poly1305_decrypt_tb_c_l60_c18_76e3_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_2_d41d_chacha20poly1305_decrypt_tb_c_l53_c25_2390_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_30_d41d_chacha20poly1305_decrypt_tb_c_l60_c27_7fac_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_31_d41d_chacha20poly1305_decrypt_tb_c_l60_c36_5acc_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_3_d41d_chacha20poly1305_decrypt_tb_c_l53_c33_c5b4_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_4_d41d_chacha20poly1305_decrypt_tb_c_l54_c9_2fa0_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_5_d41d_chacha20poly1305_decrypt_tb_c_l54_c17_ab39_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_6_d41d_chacha20poly1305_decrypt_tb_c_l54_c25_edba_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_7_d41d_chacha20poly1305_decrypt_tb_c_l54_c33_1286_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_8_d41d_chacha20poly1305_decrypt_tb_c_l55_c9_2fa1_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10 := VAR_CONST_REF_RD_uint8_t_uint8_t_32_9_d41d_chacha20poly1305_decrypt_tb_c_l55_c17_a88f_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814[chacha20poly1305_decrypt_tb_c_l42_c5_5814] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg3;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg4;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg5;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg6;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg7;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg8;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg9;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg10;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg11;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg12;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg13;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg14;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg15;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg16;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg17;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg18;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg19;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg20;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg21;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg22;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg23;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg24;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg25;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg26;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg27;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg28;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg29;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg30;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg31;
     printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l42_c5_5814_chacha20poly1305_decrypt_tb_c_l42_c5_5814_arg32;
     -- Outputs

   end if;
 end loop;

end process;

end arch;
