-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 976
entity tb_0CLK_18e0fa84 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in tb_global_to_module_t;
 module_to_global : out tb_module_to_global_t;
 return_output : out axis128_t_stream_t);
end tb_0CLK_18e0fa84;
architecture arch of tb_0CLK_18e0fa84 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal input_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal ciphertext_in_stream : uint8_t_144 := (others => to_unsigned(0, 8));
signal ciphertext_remaining_in : unsigned(31 downto 0) := to_unsigned(0, 32);
signal cycle_counter : unsigned(31 downto 0) := to_unsigned(0, 32);
signal output_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_size : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_remaining_out : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_expected : uint8_t_128 := (others => to_unsigned(0, 8));
signal tag_match_checked : unsigned(0 downto 0) := to_unsigned(0, 1);
signal chacha20poly1305_decrypt_axis_in : axis128_t_stream_t := axis128_t_stream_t_NULL;
signal REG_COMB_input_packet_count : unsigned(31 downto 0);
signal REG_COMB_ciphertext_in_stream : uint8_t_144;
signal REG_COMB_ciphertext_remaining_in : unsigned(31 downto 0);
signal REG_COMB_cycle_counter : unsigned(31 downto 0);
signal REG_COMB_output_packet_count : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_size : unsigned(31 downto 0);
signal REG_COMB_plaintext_remaining_out : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_expected : uint8_t_128;
signal REG_COMB_tag_match_checked : unsigned(0 downto 0);
signal REG_COMB_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l179_c8_7b5b]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l180_c1_7c41]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : uint8_t_144;

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : uint8_t_128;

-- printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5[chacha20poly1305_decrypt_tb_c_l181_c9_c6d5]
signal printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE : unsigned(0 downto 0);

-- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l183_c117_5672]
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x : unsigned(255 downto 0);
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output : unsigned(255 downto 0);

-- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l183_c148_a244]
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x : unsigned(255 downto 0);
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output : unsigned(255 downto 0);

-- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l183_c179_5320]
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x : unsigned(255 downto 0);
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output : unsigned(255 downto 0);

-- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l183_c210_dd6b]
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x : unsigned(255 downto 0);
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output : unsigned(255 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l183_c241_c503]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x : unsigned(255 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output : unsigned(255 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l183_c272_ff56]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x : unsigned(255 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output : unsigned(255 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l183_c302_7d05]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x : unsigned(255 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output : unsigned(255 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l183_c332_ac31]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x : unsigned(255 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output : unsigned(255 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a[chacha20poly1305_decrypt_tb_c_l183_c64_c02a]
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7 : unsigned(31 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l184_c100_991d]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x : unsigned(95 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output : unsigned(95 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l184_c130_f1af]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x : unsigned(95 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output : unsigned(95 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l184_c160_f8ee]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x : unsigned(95 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output : unsigned(95 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5[chacha20poly1305_decrypt_tb_c_l184_c65_90c5]
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2 : unsigned(31 downto 0);

-- print_aad[chacha20poly1305_decrypt_tb_c_l185_c9_cea2]
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE : unsigned(0 downto 0);
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad : uint8_t_32;
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l189_c32_b4a2]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c35_3d79]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd[chacha20poly1305_decrypt_tb_c_l191_c9_b4dd]
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l194_c30_650d]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c34_803d]
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output : uint8_t_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0[chacha20poly1305_decrypt_tb_c_l200_c9_c7e0]
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l208_c8_3bbd]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l209_c1_080f]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(31 downto 0);

-- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488]
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : axis128_t_stream_t;

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1]
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);

-- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l221_c56_fc07]
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left : unsigned(31 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right : unsigned(4 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l224_c12_5f7e]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l225_c1_fb4c]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(31 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l226_c176_f437]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l226_c207_e041]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l226_c237_7f8b]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l226_c267_c80a]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded[chacha20poly1305_decrypt_tb_c_l226_c108_8ded]
signal printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l228_c1_3d02]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c[chacha20poly1305_decrypt_tb_c_l229_c17_7c0c]
signal printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l231_c17_6e35]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l233_c17_70ec]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output : unsigned(31 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l242_c8_11d4]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_a231]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l245_c169_e848]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l245_c200_b101]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l245_c230_d9b3]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l245_c260_8481]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5[chacha20poly1305_decrypt_tb_c_l245_c105_92b5]
signal printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9]
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l262_c1_0443]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l269_c1_ae79]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l263_c16_75b7]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right : unsigned(4 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l263_c1_e17d]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l265_c1_048a]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l263_c13_e16a]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696[chacha20poly1305_decrypt_tb_c_l264_c17_0696]
signal printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68[chacha20poly1305_decrypt_tb_c_l266_c17_9a68]
signal printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0 : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l270_c16_adec]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l270_c1_917d]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da[chacha20poly1305_decrypt_tb_c_l271_c18_a6da]
signal printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l273_c17_6beb]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l280_c9_8587]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output : unsigned(0 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l280_c41_e859]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l280_c9_0d90]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l280_c69_4714]
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l280_c9_1dc0]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l281_c1_6d2f]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : uint8_t_144;

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : uint8_t_128;

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l282_c13_0ba5]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l283_c1_dfa4]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l285_c1_5a6d]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a[chacha20poly1305_decrypt_tb_c_l284_c13_746a]
signal printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0 : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f[chacha20poly1305_decrypt_tb_c_l286_c13_4b4f]
signal printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l290_c9_104d]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output : unsigned(32 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l291_c12_9b87]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l292_c1_22cd]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : uint8_t_144;

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : uint8_t_128;

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l294_c17_a7a4]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l294_c1_fccf]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : uint8_t_144;

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : uint8_t_128;

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l296_c40_e9c0]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l297_c43_4a0d]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7[chacha20poly1305_decrypt_tb_c_l298_c17_f8d7]
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l301_c38_a3f6]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l304_c42_d4b3]
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output : uint8_t_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274[chacha20poly1305_decrypt_tb_c_l306_c17_8274]
signal printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l313_c9_a764]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output : unsigned(0 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l313_c5_fec8]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l317_c5_217c]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint8_t_144_uint8_t_144_a26f( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_b938( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;

      return_output := base;
      return return_output; 
end function;

function uint8_array32_be( x : uint8_t_32) return unsigned is

  --variable x : uint8_t_32;
  variable return_output : unsigned(255 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15)&x(16)&x(17)&x(18)&x(19)&x(20)&x(21)&x(22)&x(23)&x(24)&x(25)&x(26)&x(27)&x(28)&x(29)&x(30)&x(31);
return return_output;
end function;

function uint8_array12_be( x : uint8_t_12) return unsigned is

  --variable x : uint8_t_12;
  variable return_output : unsigned(95 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11);
return return_output;
end function;

function CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_16 is
 
  variable base : axis128_t_stream_t; 
  variable return_output : uint8_t_16;
begin
      base.data.tdata(0) := ref_toks_0;
      base.data.tdata(1) := ref_toks_1;
      base.data.tdata(2) := ref_toks_2;
      base.data.tdata(3) := ref_toks_3;
      base.data.tdata(4) := ref_toks_4;
      base.data.tdata(5) := ref_toks_5;
      base.data.tdata(6) := ref_toks_6;
      base.data.tdata(7) := ref_toks_7;
      base.data.tdata(8) := ref_toks_8;
      base.data.tdata(9) := ref_toks_9;
      base.data.tdata(10) := ref_toks_10;
      base.data.tdata(11) := ref_toks_11;
      base.data.tdata(12) := ref_toks_12;
      base.data.tdata(13) := ref_toks_13;
      base.data.tdata(14) := ref_toks_14;
      base.data.tdata(15) := ref_toks_15;

      return_output := base.data.tdata;
      return return_output; 
end function;

function uint8_array16_be( x : uint8_t_16) return unsigned is

  --variable x : uint8_t_16;
  variable return_output : unsigned(127 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15);
return return_output;
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tdata(0) := ref_toks_1;
      base.data.tkeep(1) := ref_toks_2;
      base.data.tdata(1) := ref_toks_3;
      base.data.tkeep(2) := ref_toks_4;
      base.data.tdata(2) := ref_toks_5;
      base.data.tkeep(3) := ref_toks_6;
      base.data.tdata(3) := ref_toks_7;
      base.data.tkeep(4) := ref_toks_8;
      base.data.tdata(4) := ref_toks_9;
      base.data.tkeep(5) := ref_toks_10;
      base.data.tdata(5) := ref_toks_11;
      base.data.tkeep(6) := ref_toks_12;
      base.data.tdata(6) := ref_toks_13;
      base.data.tkeep(7) := ref_toks_14;
      base.data.tdata(7) := ref_toks_15;
      base.data.tkeep(8) := ref_toks_16;
      base.data.tdata(8) := ref_toks_17;
      base.data.tkeep(9) := ref_toks_18;
      base.data.tdata(9) := ref_toks_19;
      base.data.tkeep(10) := ref_toks_20;
      base.data.tdata(10) := ref_toks_21;
      base.data.tkeep(11) := ref_toks_22;
      base.data.tdata(11) := ref_toks_23;
      base.data.tkeep(12) := ref_toks_24;
      base.data.tdata(12) := ref_toks_25;
      base.data.tkeep(13) := ref_toks_26;
      base.data.tdata(13) := ref_toks_27;
      base.data.tkeep(14) := ref_toks_28;
      base.data.tdata(14) := ref_toks_29;
      base.data.tkeep(15) := ref_toks_30;
      base.data.tdata(15) := ref_toks_31;
      base.data.tlast := ref_toks_32;
      base.valid := ref_toks_33;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_32_uint8_t_32_1367( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned) return uint8_t_32 is
 
  variable base : uint8_t_32; 
  variable return_output : uint8_t_32;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;
      base(12) := ref_toks_12;
      base(13) := ref_toks_13;
      base(14) := ref_toks_14;
      base(15) := ref_toks_15;
      base(16) := ref_toks_16;
      base(17) := ref_toks_17;
      base(18) := ref_toks_18;
      base(19) := ref_toks_19;
      base(20) := ref_toks_20;
      base(21) := ref_toks_21;
      base(22) := ref_toks_22;
      base(23) := ref_toks_23;
      base(24) := ref_toks_24;
      base(25) := ref_toks_25;
      base(26) := ref_toks_26;
      base(27) := ref_toks_27;
      base(28) := ref_toks_28;
      base(29) := ref_toks_29;
      base(30) := ref_toks_30;
      base(31) := ref_toks_31;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return uint8_t_12 is
 
  variable base : uint8_t_12; 
  variable return_output : uint8_t_12;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_f92b( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned;
 ref_toks_113 : unsigned;
 ref_toks_114 : unsigned;
 ref_toks_115 : unsigned;
 ref_toks_116 : unsigned;
 ref_toks_117 : unsigned;
 ref_toks_118 : unsigned;
 ref_toks_119 : unsigned;
 ref_toks_120 : unsigned;
 ref_toks_121 : unsigned;
 ref_toks_122 : unsigned;
 ref_toks_123 : unsigned;
 ref_toks_124 : unsigned;
 ref_toks_125 : unsigned;
 ref_toks_126 : unsigned;
 ref_toks_127 : unsigned;
 ref_toks_128 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(82) := ref_toks_1;
      base(27) := ref_toks_2;
      base(91) := ref_toks_3;
      base(36) := ref_toks_4;
      base(100) := ref_toks_5;
      base(57) := ref_toks_6;
      base(2) := ref_toks_7;
      base(121) := ref_toks_8;
      base(66) := ref_toks_9;
      base(11) := ref_toks_10;
      base(75) := ref_toks_11;
      base(20) := ref_toks_12;
      base(84) := ref_toks_13;
      base(29) := ref_toks_14;
      base(93) := ref_toks_15;
      base(50) := ref_toks_16;
      base(59) := ref_toks_17;
      base(4) := ref_toks_18;
      base(123) := ref_toks_19;
      base(68) := ref_toks_20;
      base(13) := ref_toks_21;
      base(77) := ref_toks_22;
      base(22) := ref_toks_23;
      base(86) := ref_toks_24;
      base(52) := ref_toks_25;
      base(116) := ref_toks_26;
      base(61) := ref_toks_27;
      base(6) := ref_toks_28;
      base(125) := ref_toks_29;
      base(70) := ref_toks_30;
      base(15) := ref_toks_31;
      base(79) := ref_toks_32;
      base(24) := ref_toks_33;
      base(88) := ref_toks_34;
      base(45) := ref_toks_35;
      base(109) := ref_toks_36;
      base(54) := ref_toks_37;
      base(118) := ref_toks_38;
      base(63) := ref_toks_39;
      base(8) := ref_toks_40;
      base(127) := ref_toks_41;
      base(72) := ref_toks_42;
      base(17) := ref_toks_43;
      base(81) := ref_toks_44;
      base(38) := ref_toks_45;
      base(102) := ref_toks_46;
      base(47) := ref_toks_47;
      base(111) := ref_toks_48;
      base(56) := ref_toks_49;
      base(1) := ref_toks_50;
      base(120) := ref_toks_51;
      base(65) := ref_toks_52;
      base(10) := ref_toks_53;
      base(74) := ref_toks_54;
      base(31) := ref_toks_55;
      base(95) := ref_toks_56;
      base(40) := ref_toks_57;
      base(104) := ref_toks_58;
      base(49) := ref_toks_59;
      base(113) := ref_toks_60;
      base(58) := ref_toks_61;
      base(3) := ref_toks_62;
      base(122) := ref_toks_63;
      base(67) := ref_toks_64;
      base(33) := ref_toks_65;
      base(97) := ref_toks_66;
      base(42) := ref_toks_67;
      base(106) := ref_toks_68;
      base(51) := ref_toks_69;
      base(115) := ref_toks_70;
      base(60) := ref_toks_71;
      base(124) := ref_toks_72;
      base(69) := ref_toks_73;
      base(26) := ref_toks_74;
      base(90) := ref_toks_75;
      base(35) := ref_toks_76;
      base(99) := ref_toks_77;
      base(44) := ref_toks_78;
      base(108) := ref_toks_79;
      base(53) := ref_toks_80;
      base(117) := ref_toks_81;
      base(62) := ref_toks_82;
      base(126) := ref_toks_83;
      base(19) := ref_toks_84;
      base(83) := ref_toks_85;
      base(28) := ref_toks_86;
      base(92) := ref_toks_87;
      base(37) := ref_toks_88;
      base(101) := ref_toks_89;
      base(46) := ref_toks_90;
      base(110) := ref_toks_91;
      base(55) := ref_toks_92;
      base(119) := ref_toks_93;
      base(12) := ref_toks_94;
      base(76) := ref_toks_95;
      base(21) := ref_toks_96;
      base(85) := ref_toks_97;
      base(30) := ref_toks_98;
      base(94) := ref_toks_99;
      base(39) := ref_toks_100;
      base(103) := ref_toks_101;
      base(48) := ref_toks_102;
      base(112) := ref_toks_103;
      base(5) := ref_toks_104;
      base(14) := ref_toks_105;
      base(78) := ref_toks_106;
      base(23) := ref_toks_107;
      base(87) := ref_toks_108;
      base(32) := ref_toks_109;
      base(96) := ref_toks_110;
      base(41) := ref_toks_111;
      base(105) := ref_toks_112;
      base(114) := ref_toks_113;
      base(7) := ref_toks_114;
      base(71) := ref_toks_115;
      base(16) := ref_toks_116;
      base(80) := ref_toks_117;
      base(25) := ref_toks_118;
      base(89) := ref_toks_119;
      base(34) := ref_toks_120;
      base(98) := ref_toks_121;
      base(43) := ref_toks_122;
      base(107) := ref_toks_123;
      base(0) := ref_toks_124;
      base(64) := ref_toks_125;
      base(9) := ref_toks_126;
      base(73) := ref_toks_127;
      base(18) := ref_toks_128;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_128_uint8_t_128_5b48( ref_toks_0 : uint8_t_128;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned) return uint8_t_128 is
 
  variable base : uint8_t_128; 
  variable return_output : uint8_t_128;
begin
      base := ref_toks_0;
      base(108) := ref_toks_1;
      base(53) := ref_toks_2;
      base(50) := ref_toks_3;
      base(59) := ref_toks_4;
      base(4) := ref_toks_5;
      base(68) := ref_toks_6;
      base(13) := ref_toks_7;
      base(77) := ref_toks_8;
      base(10) := ref_toks_9;
      base(22) := ref_toks_10;
      base(74) := ref_toks_11;
      base(86) := ref_toks_12;
      base(19) := ref_toks_13;
      base(83) := ref_toks_14;
      base(28) := ref_toks_15;
      base(92) := ref_toks_16;
      base(37) := ref_toks_17;
      base(101) := ref_toks_18;
      base(46) := ref_toks_19;
      base(43) := ref_toks_20;
      base(110) := ref_toks_21;
      base(107) := ref_toks_22;
      base(52) := ref_toks_23;
      base(61) := ref_toks_24;
      base(6) := ref_toks_25;
      base(70) := ref_toks_26;
      base(3) := ref_toks_27;
      base(15) := ref_toks_28;
      base(79) := ref_toks_29;
      base(12) := ref_toks_30;
      base(76) := ref_toks_31;
      base(21) := ref_toks_32;
      base(85) := ref_toks_33;
      base(30) := ref_toks_34;
      base(94) := ref_toks_35;
      base(39) := ref_toks_36;
      base(36) := ref_toks_37;
      base(103) := ref_toks_38;
      base(100) := ref_toks_39;
      base(45) := ref_toks_40;
      base(109) := ref_toks_41;
      base(54) := ref_toks_42;
      base(63) := ref_toks_43;
      base(8) := ref_toks_44;
      base(72) := ref_toks_45;
      base(5) := ref_toks_46;
      base(69) := ref_toks_47;
      base(14) := ref_toks_48;
      base(78) := ref_toks_49;
      base(23) := ref_toks_50;
      base(87) := ref_toks_51;
      base(32) := ref_toks_52;
      base(29) := ref_toks_53;
      base(96) := ref_toks_54;
      base(41) := ref_toks_55;
      base(93) := ref_toks_56;
      base(38) := ref_toks_57;
      base(105) := ref_toks_58;
      base(102) := ref_toks_59;
      base(47) := ref_toks_60;
      base(111) := ref_toks_61;
      base(56) := ref_toks_62;
      base(1) := ref_toks_63;
      base(65) := ref_toks_64;
      base(62) := ref_toks_65;
      base(7) := ref_toks_66;
      base(71) := ref_toks_67;
      base(16) := ref_toks_68;
      base(80) := ref_toks_69;
      base(25) := ref_toks_70;
      base(89) := ref_toks_71;
      base(34) := ref_toks_72;
      base(31) := ref_toks_73;
      base(98) := ref_toks_74;
      base(95) := ref_toks_75;
      base(40) := ref_toks_76;
      base(104) := ref_toks_77;
      base(49) := ref_toks_78;
      base(58) := ref_toks_79;
      base(55) := ref_toks_80;
      base(67) := ref_toks_81;
      base(0) := ref_toks_82;
      base(64) := ref_toks_83;
      base(9) := ref_toks_84;
      base(73) := ref_toks_85;
      base(18) := ref_toks_86;
      base(82) := ref_toks_87;
      base(27) := ref_toks_88;
      base(24) := ref_toks_89;
      base(91) := ref_toks_90;
      base(88) := ref_toks_91;
      base(33) := ref_toks_92;
      base(97) := ref_toks_93;
      base(42) := ref_toks_94;
      base(106) := ref_toks_95;
      base(51) := ref_toks_96;
      base(48) := ref_toks_97;
      base(60) := ref_toks_98;
      base(57) := ref_toks_99;
      base(2) := ref_toks_100;
      base(66) := ref_toks_101;
      base(11) := ref_toks_102;
      base(75) := ref_toks_103;
      base(20) := ref_toks_104;
      base(17) := ref_toks_105;
      base(84) := ref_toks_106;
      base(81) := ref_toks_107;
      base(26) := ref_toks_108;
      base(90) := ref_toks_109;
      base(35) := ref_toks_110;
      base(99) := ref_toks_111;
      base(44) := ref_toks_112;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72 : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5 : entity work.printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE);

-- CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672 : 0 clocks latency
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672 : entity work.CONST_SR_224_uint256_t_0CLK_de264c78 port map (
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x,
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output);

-- CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244 : 0 clocks latency
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244 : entity work.CONST_SR_192_uint256_t_0CLK_de264c78 port map (
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x,
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output);

-- CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320 : 0 clocks latency
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320 : entity work.CONST_SR_160_uint256_t_0CLK_de264c78 port map (
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x,
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output);

-- CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b : 0 clocks latency
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b : entity work.CONST_SR_128_uint256_t_0CLK_de264c78 port map (
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x,
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503 : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503 : entity work.CONST_SR_96_uint256_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56 : entity work.CONST_SR_64_uint256_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05 : entity work.CONST_SR_32_uint256_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31 : entity work.CONST_SR_0_uint256_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a : entity work.printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d : entity work.CONST_SR_64_uint96_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af : entity work.CONST_SR_32_uint96_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee : entity work.CONST_SR_0_uint96_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5 : entity work.printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2);

-- print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2 : 0 clocks latency
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2 : entity work.print_aad_0CLK_fa355561 port map (
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE,
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad,
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2 : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2 : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd : entity work.printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0,
printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d : 0 clocks latency
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d : entity work.VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0 : entity work.printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0,
printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : 0 clocks latency
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488 : entity work.MUX_uint1_t_axis128_t_stream_t_axis128_t_stream_t_0CLK_de264c78 port map (
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

-- BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07 : 0 clocks latency
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07 : entity work.BIN_OP_LTE_uint32_t_uint5_t_0CLK_e595f783 port map (
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437 : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437 : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded : entity work.printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0,
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1,
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2,
printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c : entity work.printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848 : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848 : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481 : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5 : entity work.printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0,
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1,
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2,
printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7 : entity work.BIN_OP_GT_uint32_t_uint5_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696 : entity work.printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE);

-- printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68 : entity work.printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da : entity work.printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output);

-- UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714 : 0 clocks latency
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr,
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52 : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5 : entity work.BIN_OP_EQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a : entity work.printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0);

-- printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f : entity work.printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854 : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4 : entity work.BIN_OP_EQ_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5 : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0 : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0 : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7 : entity work.printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0,
printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3 : 0 clocks latency
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3 : entity work.VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274 : entity work.printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0,
printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764 : entity work.BIN_OP_GT_uint32_t_uint32_t_0CLK_380ecc95 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a : 0 clocks latency
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a : entity work.BIN_OP_MINUS_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 input_packet_count,
 ciphertext_in_stream,
 ciphertext_remaining_in,
 cycle_counter,
 output_packet_count,
 plaintext_out_size,
 plaintext_remaining_out,
 plaintext_out_expected,
 tag_match_checked,
 chacha20poly1305_decrypt_axis_in,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
 CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output,
 CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output,
 CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output,
 CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output,
 VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
 BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output,
 UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output,
 VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output,
 BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_key : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_nonce : uint8_t_12;
 variable VAR_chacha20poly1305_decrypt_aad : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_aad_len : unsigned(7 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_tags_match : unsigned(0 downto 0);
 variable VAR_key : uint8_t_32;
 variable VAR_nonce : uint8_t_12;
 variable VAR_aad : uint8_t_32;
 variable VAR_aad_len : unsigned(31 downto 0);
 variable VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_f60f_0 : unsigned(31 downto 0);
 variable VAR_plaintexts : uint8_t_2_128;
 variable VAR_plaintext_lens : uint32_t_2;
 variable VAR_input_ciphertext0 : uint8_t_144;
 variable VAR_input_ciphertext1 : uint8_t_144;
 variable VAR_input_ciphertexts : uint8_t_2_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_2261_return_output : uint8_t_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_1997_return_output : uint8_t_144;
 variable VAR_ciphertext_lens : uint32_t_2;
 variable VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_f10d : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_6f9e : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_84c1 : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_PRINT_32_BYTES_uint : unsigned(255 downto 0);
 variable VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x : unsigned(255 downto 0);
 variable VAR_PRINT_12_BYTES_uint : unsigned(95 downto 0);
 variable VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_7d68_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x : unsigned(95 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad : uint8_t_32;
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len : unsigned(31 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output : uint8_t_array_128_t;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0 : uint8_t_128;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1 : uint8_t_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond : unsigned(0 downto 0);
 variable VAR_i : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond : unsigned(0 downto 0);
 variable VAR_PRINT_16_BYTES_uint : unsigned(127 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l226_c62_8b02_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x : unsigned(127 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l231_c17_66ef : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output : unsigned(31 downto 0);
 variable VAR_ARRAY_SHIFT_DOWN_i : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l242_c8_9478_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l245_c58_481d_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x : unsigned(127 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_pos : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l296_c17_3517 : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l304_c17_0020 : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output : uint8_t_array_128_t;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0 : uint8_t_128;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1 : uint8_t_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond : unsigned(0 downto 0);
 variable VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l317_c5_30ca : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l158_l183_DUPLICATE_45c3_return_output : uint8_t_32;
 variable VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_01f5_return_output : uint8_t_12;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_4a53_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9326_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_6f11_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f6fa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f368_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_44ed_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_8570_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0dbc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_1fca_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_3d4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_a444_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9b24_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_6c44_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_c57d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_4b3e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0356_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a_return_output : uint8_t_144;
 variable VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a_return_output : uint8_t_128;
 -- State registers comb logic variables
variable REG_VAR_input_packet_count : unsigned(31 downto 0);
variable REG_VAR_ciphertext_in_stream : uint8_t_144;
variable REG_VAR_ciphertext_remaining_in : unsigned(31 downto 0);
variable REG_VAR_cycle_counter : unsigned(31 downto 0);
variable REG_VAR_output_packet_count : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_size : unsigned(31 downto 0);
variable REG_VAR_plaintext_remaining_out : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_expected : uint8_t_128;
variable REG_VAR_tag_match_checked : unsigned(0 downto 0);
variable REG_VAR_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_input_packet_count := input_packet_count;
  REG_VAR_ciphertext_in_stream := ciphertext_in_stream;
  REG_VAR_ciphertext_remaining_in := ciphertext_remaining_in;
  REG_VAR_cycle_counter := cycle_counter;
  REG_VAR_output_packet_count := output_packet_count;
  REG_VAR_plaintext_out_size := plaintext_out_size;
  REG_VAR_plaintext_remaining_out := plaintext_remaining_out;
  REG_VAR_plaintext_out_expected := plaintext_out_expected;
  REG_VAR_tag_match_checked := tag_match_checked;
  REG_VAR_chacha20poly1305_decrypt_axis_in := chacha20poly1305_decrypt_axis_in;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(1, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue := to_unsigned(0, 1);
     VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_f60f_0 := to_unsigned(29, 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len := VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_f60f_0;
     VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_f10d := resize(VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_f60f_0, 8);
     VAR_chacha20poly1305_decrypt_aad_len := VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_f10d;
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(14, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(15, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right := to_unsigned(1, 1);
     VAR_chacha20poly1305_decrypt_axis_out_ready := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(4, 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad := to_byte_array("Additional authenticated data", 32);
     VAR_chacha20poly1305_decrypt_aad := to_byte_array("Additional authenticated data", 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(3, 32);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(6, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(5, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(9, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1 := to_unsigned(71, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1 := to_unsigned(71, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right := to_unsigned(0, 1);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue := to_unsigned(0, 1);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := to_unsigned(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(11, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(7, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left := to_unsigned(0, 1);
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right := to_unsigned(16, 5);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse := to_unsigned(0, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0 := to_unsigned(80, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0 := to_unsigned(80, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse := to_unsigned(0, 8);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(15, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(15, 32);
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse := to_unsigned(0, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(8, 32);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(5, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0 := to_unsigned(56, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0 := to_unsigned(56, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(3, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(10, 32);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right := to_unsigned(2, 2);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1 := to_unsigned(96, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1 := to_unsigned(96, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(8, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right := to_signed(0, 32);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right := to_unsigned(16, 5);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right := to_signed(12, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse := to_unsigned(0, 1);
     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l282_c13_0ba5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output;

     -- CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l158_l183_DUPLICATE_45c3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l158_l183_DUPLICATE_45c3_return_output := CONST_REF_RD_uint8_t_32_uint8_t_32_1367(
     to_unsigned(128, 8),
     to_unsigned(129, 8),
     to_unsigned(130, 8),
     to_unsigned(131, 8),
     to_unsigned(132, 8),
     to_unsigned(133, 8),
     to_unsigned(134, 8),
     to_unsigned(135, 8),
     to_unsigned(136, 8),
     to_unsigned(137, 8),
     to_unsigned(138, 8),
     to_unsigned(139, 8),
     to_unsigned(140, 8),
     to_unsigned(141, 8),
     to_unsigned(142, 8),
     to_unsigned(143, 8),
     to_unsigned(144, 8),
     to_unsigned(145, 8),
     to_unsigned(146, 8),
     to_unsigned(147, 8),
     to_unsigned(148, 8),
     to_unsigned(149, 8),
     to_unsigned(150, 8),
     to_unsigned(151, 8),
     to_unsigned(152, 8),
     to_unsigned(153, 8),
     to_unsigned(154, 8),
     to_unsigned(155, 8),
     to_unsigned(156, 8),
     to_unsigned(157, 8),
     to_unsigned(158, 8),
     to_unsigned(159, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_b938[chacha20poly1305_decrypt_tb_c_l150_c9_1997] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_1997_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_b938(
     (others => to_unsigned(0, 8)),
     to_unsigned(207, 8),
     to_unsigned(18, 8),
     to_unsigned(153, 8),
     to_unsigned(56, 8),
     to_unsigned(109, 8),
     to_unsigned(148, 8),
     to_unsigned(46, 8),
     to_unsigned(223, 8),
     to_unsigned(86, 8),
     to_unsigned(194, 8),
     to_unsigned(230, 8),
     to_unsigned(136, 8),
     to_unsigned(22, 8),
     to_unsigned(245, 8),
     to_unsigned(98, 8),
     to_unsigned(203, 8),
     to_unsigned(225, 8),
     to_unsigned(162, 8),
     to_unsigned(237, 8),
     to_unsigned(76, 8),
     to_unsigned(125, 8),
     to_unsigned(33, 8),
     to_unsigned(38, 8),
     to_unsigned(154, 8),
     to_unsigned(145, 8),
     to_unsigned(170, 8),
     to_unsigned(177, 8),
     to_unsigned(245, 8),
     to_unsigned(58, 8),
     to_unsigned(247, 8),
     to_unsigned(109, 8),
     to_unsigned(193, 8),
     to_unsigned(110, 8),
     to_unsigned(164, 8),
     to_unsigned(226, 8),
     to_unsigned(24, 8),
     to_unsigned(224, 8),
     to_unsigned(235, 8),
     to_unsigned(42, 8),
     to_unsigned(12, 8),
     to_unsigned(203, 8),
     to_unsigned(250, 8),
     to_unsigned(213, 8),
     to_unsigned(96, 8),
     to_unsigned(218, 8),
     to_unsigned(152, 8),
     to_unsigned(26, 8),
     to_unsigned(161, 8),
     to_unsigned(57, 8),
     to_unsigned(77, 8),
     to_unsigned(241, 8),
     to_unsigned(6, 8),
     to_unsigned(215, 8),
     to_unsigned(25, 8),
     to_unsigned(30, 8),
     to_unsigned(111, 8),
     to_unsigned(55, 8),
     to_unsigned(205, 8),
     to_unsigned(247, 8),
     to_unsigned(170, 8),
     to_unsigned(118, 8),
     to_unsigned(205, 8),
     to_unsigned(122, 8),
     to_unsigned(43, 8),
     to_unsigned(152, 8),
     to_unsigned(145, 8),
     to_unsigned(176, 8),
     to_unsigned(58, 8),
     to_unsigned(35, 8),
     to_unsigned(116, 8),
     to_unsigned(207, 8),
     to_unsigned(172, 8),
     to_unsigned(236, 8),
     to_unsigned(106, 8),
     to_unsigned(222, 8),
     to_unsigned(195, 8),
     to_unsigned(78, 8),
     to_unsigned(102, 8),
     to_unsigned(105, 8),
     to_unsigned(120, 8),
     to_unsigned(7, 8),
     to_unsigned(199, 8),
     to_unsigned(227, 8),
     to_unsigned(31, 8),
     to_unsigned(15, 8),
     to_unsigned(235, 8),
     to_unsigned(75, 8),
     to_unsigned(97, 8),
     to_unsigned(234, 8),
     to_unsigned(45, 8),
     to_unsigned(210, 8),
     to_unsigned(164, 8),
     to_unsigned(89, 8),
     to_unsigned(124, 8),
     to_unsigned(174, 8),
     to_unsigned(233, 8));

     -- CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_01f5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_01f5_return_output := CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2(
     to_unsigned(7, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(64, 8),
     to_unsigned(65, 8),
     to_unsigned(66, 8),
     to_unsigned(67, 8),
     to_unsigned(68, 8),
     to_unsigned(69, 8),
     to_unsigned(70, 8),
     to_unsigned(71, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_a26f[chacha20poly1305_decrypt_tb_c_l149_c9_2261] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_2261_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_a26f(
     (others => to_unsigned(0, 8)),
     to_unsigned(215, 8),
     to_unsigned(30, 8),
     to_unsigned(133, 8),
     to_unsigned(49, 8),
     to_unsigned(110, 8),
     to_unsigned(221, 8),
     to_unsigned(3, 8),
     to_unsigned(242, 8),
     to_unsigned(92, 8),
     to_unsigned(174, 8),
     to_unsigned(198, 8),
     to_unsigned(184, 8),
     to_unsigned(94, 8),
     to_unsigned(232, 8),
     to_unsigned(122, 8),
     to_unsigned(221, 8),
     to_unsigned(225, 8),
     to_unsigned(237, 8),
     to_unsigned(168, 8),
     to_unsigned(104, 8),
     to_unsigned(96, 8),
     to_unsigned(115, 8),
     to_unsigned(11, 8),
     to_unsigned(185, 8),
     to_unsigned(168, 8),
     to_unsigned(235, 8),
     to_unsigned(162, 8),
     to_unsigned(227, 8),
     to_unsigned(117, 8),
     to_unsigned(246, 8),
     to_unsigned(102, 8),
     to_unsigned(196, 8),
     to_unsigned(35, 8),
     to_unsigned(178, 8),
     to_unsigned(235, 8),
     to_unsigned(84, 8),
     to_unsigned(201, 8),
     to_unsigned(250, 8),
     to_unsigned(121, 8),
     to_unsigned(88, 8),
     to_unsigned(152, 8),
     to_unsigned(174, 8),
     to_unsigned(215, 8),
     to_unsigned(124, 8),
     to_unsigned(142, 8),
     to_unsigned(251, 8),
     to_unsigned(38, 8),
     to_unsigned(128, 8),
     to_unsigned(28, 8),
     to_unsigned(119, 8),
     to_unsigned(146, 8),
     to_unsigned(15, 8),
     to_unsigned(219, 8),
     to_unsigned(8, 8),
     to_unsigned(9, 8),
     to_unsigned(110, 8),
     to_unsigned(96, 8),
     to_unsigned(164, 8),
     to_unsigned(133, 8),
     to_unsigned(207, 8),
     to_unsigned(17, 8),
     to_unsigned(184, 8),
     to_unsigned(27, 8),
     to_unsigned(89, 8),
     to_unsigned(93, 8),
     to_unsigned(168, 8),
     to_unsigned(125, 8),
     to_unsigned(106, 8),
     to_unsigned(45, 8),
     to_unsigned(3, 8),
     to_unsigned(201, 8),
     to_unsigned(186, 8),
     to_unsigned(223, 8),
     to_unsigned(92, 8),
     to_unsigned(185, 8),
     to_unsigned(71, 8),
     to_unsigned(116, 8),
     to_unsigned(66, 8),
     to_unsigned(18, 8),
     to_unsigned(63, 8));

     -- Submodule level 1
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_1997_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_1997_return_output;
     VAR_chacha20poly1305_decrypt_key := VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l158_l183_DUPLICATE_45c3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l282_c13_0ba5_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_2261_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_2261_return_output;
     VAR_chacha20poly1305_decrypt_nonce := VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_01f5_return_output;
     -- uint8_array32_be[chacha20poly1305_decrypt_tb_c_l183_c41_2dde] LATENCY=0
     VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output := uint8_array32_be(
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l158_l183_DUPLICATE_45c3_return_output);

     -- uint8_array12_be[chacha20poly1305_decrypt_tb_c_l184_c40_7d68] LATENCY=0
     VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_7d68_return_output := uint8_array12_be(
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_01f5_return_output);

     -- Submodule level 2
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_7d68_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_7d68_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_7d68_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_2dde_return_output;
     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l183_c302_7d05] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output;

     -- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l183_c179_5320] LATENCY=0
     -- Inputs
     CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x <= VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_x;
     -- Outputs
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output := CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l183_c272_ff56] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l184_c160_f8ee] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l184_c100_991d] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l183_c241_c503] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output;

     -- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l183_c210_dd6b] LATENCY=0
     -- Inputs
     CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x <= VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_x;
     -- Outputs
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output := CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l184_c130_f1af] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l183_c332_ac31] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output;

     -- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l183_c148_a244] LATENCY=0
     -- Inputs
     CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x <= VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_x;
     -- Outputs
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output := CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output;

     -- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l183_c117_5672] LATENCY=0
     -- Inputs
     CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x <= VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_x;
     -- Outputs
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output := CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1 := resize(VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_a244_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3 := resize(VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_dd6b_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_f8ee_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_c503_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2 := resize(VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_5320_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_ac31_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_f1af_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_7d05_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_ff56_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0 := resize(VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_5672_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_991d_return_output, 32);
 -- Reads from global variables
     VAR_chacha20poly1305_decrypt_axis_in_ready := global_to_module.chacha20poly1305_decrypt_axis_in_ready;
     VAR_chacha20poly1305_decrypt_axis_out := global_to_module.chacha20poly1305_decrypt_axis_out;
     -- Submodule level 0
     VAR_return_output := VAR_chacha20poly1305_decrypt_axis_out;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right := VAR_chacha20poly1305_decrypt_axis_in_ready;
     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d[chacha20poly1305_decrypt_tb_c_l245_c58_481d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l245_c58_481d_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f368 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f368_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(4);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_6f11 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_6f11_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(2);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_44ed LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_44ed_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(5);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d[chacha20poly1305_decrypt_tb_c_l242_c8_9478] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l242_c8_9478_return_output := VAR_chacha20poly1305_decrypt_axis_out.valid;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9326 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9326_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(1);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_a444 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_a444_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(10);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f6fa LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f6fa_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(3);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_3d4b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_3d4b_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(9);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9b24 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9b24_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(11);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d[chacha20poly1305_decrypt_tb_c_l262_c12_2280] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tlast;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0356 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0356_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(15);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_1fca LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_1fca_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(8);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_4a53 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_4a53_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(0);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_4b3e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_4b3e_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(14);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0dbc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0dbc_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(7);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_8570 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_8570_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(6);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_c57d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_c57d_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(13);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_6c44 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_6c44_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(12);

     -- Submodule level 1
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_4b3e_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_4b3e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9b24_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9b24_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l262_c12_2280_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f368_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f368_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_44ed_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_44ed_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_1fca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_1fca_return_output, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l242_c8_9478_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f6fa_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_f6fa_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0dbc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0dbc_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_3d4b_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_3d4b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_4a53_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_4a53_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_a444_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_a444_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_6f11_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_6f11_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_6c44_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l252_l256_DUPLICATE_6c44_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0356_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_0356_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_c57d_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_c57d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9326_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_9326_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_8570_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l252_DUPLICATE_8570_return_output;
     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l245_c41_641a] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l245_c58_481d_return_output);

     -- Submodule level 2
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l245_c41_641a_return_output;
     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l245_c230_d9b3] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l245_c260_8481] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l245_c200_b101] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l245_c169_e848] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l245_c260_8481_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l245_c200_b101_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l245_c230_d9b3_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l245_c169_e848_return_output, 32);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue := VAR_CLOCK_ENABLE;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := ciphertext_in_stream;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := ciphertext_remaining_in;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left := input_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0 := resize(input_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0 := resize(input_packet_count, 1);
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0 := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0 := input_packet_count;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left := output_packet_count;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left := output_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0 := resize(output_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0 := resize(output_packet_count, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0 := output_packet_count;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := plaintext_out_expected;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := plaintext_out_size;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := plaintext_remaining_out;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse := tag_match_checked;
     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l242_c8_11d4] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;

     -- chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee(
     chacha20poly1305_decrypt_axis_in,
     to_unsigned(0, 1));

     -- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c34_803d] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_0;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_ref_toks_1;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output := VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l280_c41_e859] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l179_c8_7b5b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c35_3d79] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l290_c9_104d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output;

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l189_c32_b4a2] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l224_c12_5f7e] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l317_c5_217c] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l231_c17_6e35] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l194_c30_650d] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l224_c12_5f7e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l242_c8_11d4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_7b5b_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l280_c41_e859_return_output;
     VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l231_c17_66ef := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l231_c17_6e35_return_output, 32);
     VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l290_c9_104d_return_output, 32);
     VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l317_c5_30ca := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l317_c5_217c_return_output, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_3d79_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_650d_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_84c1 := VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_803d_return_output.data;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_6f9e := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_b4a2_return_output.data;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_6f9e;
     REG_VAR_cycle_counter := VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l317_c5_30ca;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l231_c17_66ef;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f, 1);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0 := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l290_c9_295f;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_84c1;
     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l180_c1_7c41] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l301_c38_a3f6] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_a231] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l304_c42_d4b3] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_0;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_ref_toks_1;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output := VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_ae72] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l291_c12_9b87] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;

     -- Submodule level 2
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l291_c12_9b87_return_output;
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7c41_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_a231_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l301_c38_a3f6_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l304_c17_0020 := VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l304_c42_d4b3_return_output.data;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output, 33)));
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l304_c17_0020;
     -- CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(10);

     -- printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5[chacha20poly1305_decrypt_tb_c_l245_c105_92b5] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_chacha20poly1305_decrypt_tb_c_l245_c105_92b5_arg3;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(41);

     -- CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(19);

     -- CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(91);

     -- CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(20);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(105);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(124);

     -- CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(59);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(37);

     -- CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(47);

     -- CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(31);

     -- CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(60);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(78);

     -- CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(74);

     -- CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(37);

     -- CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(78);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(135);

     -- CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(10);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(104);

     -- CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(50);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l208_c8_3bbd] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(1);

     -- CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(81);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(97);

     -- CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(39);

     -- CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(40);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(140);

     -- CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(101);

     -- CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(33);

     -- CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(116);

     -- CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(104);

     -- CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(55);

     -- CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(54);

     -- CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(67);

     -- CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(2);

     -- CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(38);

     -- CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(49);

     -- CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(12);

     -- CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(72);

     -- CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(93);

     -- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l221_c56_fc07] LATENCY=0
     -- Inputs
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_left;
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_right;
     -- Outputs
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output := BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(50);

     -- CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(0);

     -- CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(69);

     -- CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(61);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(16);

     -- CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(21);

     -- CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(65);

     -- CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(52);

     -- CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(56);

     -- CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(30);

     -- CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(8);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(116);

     -- CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(84);

     -- CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(100);

     -- CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(70);

     -- CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(15);

     -- CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(24);

     -- CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(109);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(139);

     -- CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(80);

     -- CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(19);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(132);

     -- CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(105);

     -- CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(93);

     -- CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(23);

     -- CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(5);

     -- CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(26);

     -- CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(32);

     -- CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(99);

     -- CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(56);

     -- CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(43);

     -- CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(82);

     -- CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(53);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(121);

     -- CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(46);

     -- CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(24);

     -- CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(28);

     -- CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(107);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(22);

     -- CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(46);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(138);

     -- CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(65);

     -- CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(71);

     -- printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5[chacha20poly1305_decrypt_tb_c_l184_c65_90c5] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_chacha20poly1305_decrypt_tb_c_l184_c65_90c5_arg2;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(52);

     -- CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(72);

     -- CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(74);

     -- CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(21);

     -- CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(8);

     -- CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(103);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(117);

     -- CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(110);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(125);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(57);

     -- CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(57);

     -- CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(44);

     -- CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(110);

     -- CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(64);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(44);

     -- CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(82);

     -- CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(85);

     -- CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(36);

     -- CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(94);

     -- CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(103);

     -- CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(34);

     -- CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(23);

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l269_c1_ae79] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(92);

     -- CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(95);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(4);

     -- CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(33);

     -- CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(30);

     -- CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(48);

     -- CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(73);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(99);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(15);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(118);

     -- CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(63);

     -- CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(25);

     -- CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(63);

     -- CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(92);

     -- CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(107);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(127);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(126);

     -- CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(115);

     -- CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(42);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(53);

     -- CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(120);

     -- CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(6);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(142);

     -- CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(95);

     -- CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(77);

     -- CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(124);

     -- CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(125);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(130);

     -- CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(81);

     -- CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(89);

     -- CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(83);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(115);

     -- CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(17);

     -- CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(58);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l233_c17_70ec] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(111);

     -- CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(45);

     -- CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(109);

     -- CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(32);

     -- printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0[chacha20poly1305_decrypt_tb_c_l200_c9_c7e0] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_chacha20poly1305_decrypt_tb_c_l200_c9_c7e0_arg1;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(83);

     -- CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(29);

     -- CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(51);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(117);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(143);

     -- CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(84);

     -- CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(17);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(126);

     -- CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(11);

     -- printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a[chacha20poly1305_decrypt_tb_c_l183_c64_c02a] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg3;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg4;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg5;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg6;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_chacha20poly1305_decrypt_tb_c_l183_c64_c02a_arg7;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(7);

     -- CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(66);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(59);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(106);

     -- CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(66);

     -- CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(97);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(89);

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l270_c16_adec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(73);

     -- CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(62);

     -- CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(100);

     -- CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(18);

     -- CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(62);

     -- CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(85);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(122);

     -- CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(25);

     -- CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(28);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(133);

     -- CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(7);

     -- CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(61);

     -- CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(11);

     -- CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(88);

     -- CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(47);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(14);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(128);

     -- CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(26);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(120);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(35);

     -- CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(102);

     -- CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(5);

     -- CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(79);

     -- CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(90);

     -- CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(69);

     -- CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(29);

     -- CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(9);

     -- CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(4);

     -- CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(27);

     -- CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(64);

     -- CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(102);

     -- CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(121);

     -- CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(60);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(141);

     -- CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(38);

     -- CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(96);

     -- CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(51);

     -- CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(18);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l280_c69_4714] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr <= VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output := UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(58);

     -- CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(2);

     -- CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(43);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(79);

     -- CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(68);

     -- CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(118);

     -- CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(80);

     -- CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(12);

     -- print_aad[chacha20poly1305_decrypt_tb_c_l185_c9_cea2] LATENCY=0
     -- Clock enable
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_CLOCK_ENABLE;
     -- Inputs
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad;
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_cea2_aad_len;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd[chacha20poly1305_decrypt_tb_c_l191_c9_b4dd] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_chacha20poly1305_decrypt_tb_c_l191_c9_b4dd_arg1;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(86);

     -- CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(40);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l263_c16_75b7] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(119);

     -- CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(127);

     -- CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(87);

     -- CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(31);

     -- printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5[chacha20poly1305_decrypt_tb_c_l181_c9_c6d5] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_chacha20poly1305_decrypt_tb_c_l181_c9_c6d5_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(14);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(136);

     -- CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(98);

     -- CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(27);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(113);

     -- CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(106);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(137);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(1);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(134);

     -- CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(55);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(90);

     -- CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(86);

     -- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_left;
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output := BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(96);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(129);

     -- CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(77);

     -- CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(9);

     -- CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(36);

     -- CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(98);

     -- CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(71);

     -- CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(75);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l273_c17_6beb] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(22);

     -- CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(111);

     -- CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(20);

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l250_c16_e416] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(3);

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l262_c1_0443] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(16);

     -- CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(45);

     -- CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(101);

     -- CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(94);

     -- CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(0);

     -- CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(113);

     -- CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(39);

     -- CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(34);

     -- CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(6);

     -- CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(48);

     -- CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(42);

     -- CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(54);

     -- CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(49);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(70);

     -- CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(87);

     -- CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(68);

     -- FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d[chacha20poly1305_decrypt_tb_c_l274_c168_2060] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(119);

     -- CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(122);

     -- CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(75);

     -- CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(91);

     -- CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(3);

     -- CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(41);

     -- CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(35);

     -- CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(88);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d[chacha20poly1305_decrypt_tb_c_l234_c173_465e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output(131);

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l215_c16_7675] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_left;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l270_c16_adec_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l208_c8_3bbd_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l263_c16_75b7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l233_c17_70ec_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l273_c17_6beb_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l254_DUPLICATE_057a_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output, 32);
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l256_l252_DUPLICATE_5d1b_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_e257_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_403f_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_1f79_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_5f37_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l262_l242_DUPLICATE_0c81_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_4976_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3bbf_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_304b_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_fb43_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_2505_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output, 32);
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_68a7_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_dca2_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_a291_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output, 32);
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_8191_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output, 32);
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_58d3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output, 32);
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_9b06_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output, 32);
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l270_l252_DUPLICATE_0b34_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output, 32);
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l252_l270_l256_l242_DUPLICATE_a711_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_338f_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5351_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_4ed8_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_220c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output, 32);
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_3cdf_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_a13e_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_2044_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_6713_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_d108_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_3da6_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_2a91_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_6eae_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l242_l270_DUPLICATE_e3c8_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7606_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_4b62_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output, 32);
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l256_l252_l270_DUPLICATE_18ec_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ea29_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_1fc3_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_072c_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5045_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_af4f_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1b9e_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7b17_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5cff_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_fbb1_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_9093_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output, 32);
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l252_l270_l242_l256_l262_DUPLICATE_4837_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_b4c7_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_848d_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_5091_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_4c73_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_b8a9_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_6584_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l270_l274_DUPLICATE_700f_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l274_l242_DUPLICATE_fa4e_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_929e_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e076_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output, 32);
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_da86_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_306b_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l274_l242_l262_l270_DUPLICATE_e79d_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_7438_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_65d8_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_bd50_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_4dc6_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_70c5_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_e4c7_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l242_l270_l274_l262_DUPLICATE_4d7f_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_5f8e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output, 32);
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l270_l256_l242_l262_l252_DUPLICATE_dfa8_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_b4f0_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_cf22_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_b667_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_7e61_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_50a2_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_8ce4_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_961b_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1fe5_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1ed1_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_3e75_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output, 32);
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_3c30_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_2a31_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_bd6e_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_472d_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c1a5_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l262_l242_l270_l274_DUPLICATE_e947_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l274_l270_l242_l262_DUPLICATE_cbd5_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f233_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_e90f_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_4528_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_94a1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output, 32);
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_e45b_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_c762_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_3b16_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_0a89_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_68d2_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l270_l274_l242_l262_DUPLICATE_3ae6_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l270_l242_l274_DUPLICATE_d37f_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d024_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_f226_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_d0ea_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_f57f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output, 32);
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l270_l252_l242_l262_l256_DUPLICATE_6854_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_c7bb_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ba8a_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l242_l274_l262_l270_DUPLICATE_c5de_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l242_l262_l274_l270_DUPLICATE_0f96_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_1508_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l274_l262_l270_l242_DUPLICATE_e693_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l262_l274_l270_l242_DUPLICATE_c9f1_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_21f5_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l262_l274_DUPLICATE_ab9c_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l270_l242_l274_l262_DUPLICATE_ca1c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output, 32);
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l256_l270_l242_l252_l262_DUPLICATE_d334_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_f98c_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1c92_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_975b_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_d1af_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_44f7_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_ffd4_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6937_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_d33a_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_36b1_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_9811_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_831f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_6b79_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_7694_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_55e3_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_b276_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_b726_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_766a_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_ad3a_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_7b08_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_f8cb_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_ce8c_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_3b94_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_8d37_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_dfc6_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_0a5a_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_285f_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_82df_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_ea21_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_2180_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_61ea_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_dd5b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l208_l224_DUPLICATE_5426_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l208_l217_l228_l224_DUPLICATE_9cdb_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_17f3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_6905_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_9b86_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_0dd1_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_83ce_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_6562_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_c99e_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_1397_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_983d_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_a92a_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_706a_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_2655_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_708d_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_ac0a_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_f3d4_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_8046_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_c5e4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l217_l208_DUPLICATE_072c_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_232f_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_3742_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f34c_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_061c_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_8080_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l228_l234_DUPLICATE_8e0e_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_5471_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_7c67_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_f548_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_88ee_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l217_l228_DUPLICATE_a65b_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7a6_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_8f11_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_9828_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_295c_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6dea_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_8a0d_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_ccfd_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_37c6_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l208_l224_DUPLICATE_5136_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5453_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l228_l217_l224_l208_DUPLICATE_ffec_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_50db_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_8448_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_0625_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_f9b7_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_85de_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_a9c9_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_f7d5_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_e929_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_eddb_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l234_DUPLICATE_6b2b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l217_l224_DUPLICATE_a905_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l208_l224_DUPLICATE_6203_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_bddc_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_830f_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_5718_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l228_l224_DUPLICATE_7653_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l208_l224_l234_l228_DUPLICATE_2195_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_d391_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l208_l234_DUPLICATE_646b_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_bfbe_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l208_l228_DUPLICATE_66a6_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l217_l224_l208_l228_DUPLICATE_1e51_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_5eb3_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_6ca8_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l234_l208_DUPLICATE_63d6_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_4307_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_e84e_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_a408_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_7bd5_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_20df_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_511c_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_acc0_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l217_l228_l224_l208_DUPLICATE_2ae0_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_75fd_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_b154_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_2f8b_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l234_DUPLICATE_bdc1_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l208_l234_l228_l224_DUPLICATE_26b5_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l234_l208_l224_l228_DUPLICATE_1829_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l234_l228_DUPLICATE_4dd9_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_25bd_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_0d1b_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l234_l224_l228_l208_DUPLICATE_492e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l224_l217_DUPLICATE_b615_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l224_l228_l234_l208_DUPLICATE_295e_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l224_l208_l228_l234_DUPLICATE_c266_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l228_l208_DUPLICATE_4c7c_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l234_l228_l224_l208_DUPLICATE_fcff_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l234_l224_DUPLICATE_fe86_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_afc1_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l228_l234_l224_l208_DUPLICATE_167c_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l208_l228_l234_l224_DUPLICATE_1ea4_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l224_l234_l208_l228_DUPLICATE_62c0_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l228_l208_l224_l234_DUPLICATE_56f2_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l228_l224_l208_l217_DUPLICATE_1170_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_ae79_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l215_c16_7675_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c46_650b_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l234_c173_465e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l250_c16_e416_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l274_c46_3763_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l274_c168_2060_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_0443_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right := VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l280_c69_4714_return_output;
     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l265_c1_048a] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l263_c13_e16a] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l270_c1_917d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l263_c1_e17d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l209_c1_080f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l251_c1_9c01] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l252_c20_ef14] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l228_c13_5633] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l270_c13_0431] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l254_c47_6da9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l215_c13_01f1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output;

     -- Submodule level 4
     VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l265_c1_048a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l252_c20_ef14_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l254_c47_6da9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l251_c1_9c01_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l209_c1_080f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l263_c1_e17d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l270_c1_917d_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c13_5633_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l263_c13_e16a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l270_c13_0431_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l254_c30_59b7_0;
     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c(
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l221_c56_fc07_return_output,
     to_unsigned(1, 1));

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696[chacha20poly1305_decrypt_tb_c_l264_c17_0696] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l264_c17_0696_chacha20poly1305_decrypt_tb_c_l264_c17_0696_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68[chacha20poly1305_decrypt_tb_c_l266_c17_9a68] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_chacha20poly1305_decrypt_tb_c_l266_c17_9a68_arg0;
     -- Outputs

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da[chacha20poly1305_decrypt_tb_c_l271_c18_a6da] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_chacha20poly1305_decrypt_tb_c_l271_c18_a6da_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed[chacha20poly1305_decrypt_tb_c_l226_c62_8b02] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l226_c62_8b02_return_output := CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed(
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l211_c9_87a8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l215_c13_01f1_return_output);

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l225_c1_fb4c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l224_c9_1b2b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_6117] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output := FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l262_c9_aea7] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;

     -- Submodule level 5
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_6117_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l225_c1_fb4c_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l224_c9_1b2b_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c9_aea7_return_output;
     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l226_c45_f860] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l226_c62_8b02_return_output);

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l228_c1_3d02] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9[chacha20poly1305_decrypt_tb_c_l255_c21_edb9] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l248_c9_5b54_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_chacha20poly1305_decrypt_tb_c_l255_c21_edb9_arg2;
     -- Outputs

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l242_c5_8bbd] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l208_c5_d488] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;

     -- Submodule level 6
     VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l228_c1_3d02_return_output;
     REG_VAR_chacha20poly1305_decrypt_axis_in := VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output, 1);
     REG_VAR_input_packet_count := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0 := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l226_c45_f860_return_output;
     -- CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_f92b(
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output,
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l208_c5_d488_return_output);

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l280_c9_8587] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l226_c267_c80a] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l294_c17_a7a4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;

     -- CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a_return_output := CONST_REF_RD_uint8_t_128_uint8_t_128_5b48(
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_ae72_return_output,
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output,
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l242_c5_8bbd_return_output);

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l297_c43_4a0d] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l226_c207_e041] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l226_c237_7f8b] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output;

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l296_c40_e9c0] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c[chacha20poly1305_decrypt_tb_c_l229_c17_7c0c] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_chacha20poly1305_decrypt_tb_c_l229_c17_7c0c_arg0;
     -- Outputs

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l226_c176_f437] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output;

     -- Submodule level 7
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l280_c9_8587_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l294_c17_a7a4_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_5b48_chacha20poly1305_decrypt_tb_c_l280_l294_l291_DUPLICATE_130a_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_f92b_chacha20poly1305_decrypt_tb_c_l291_l280_l294_DUPLICATE_214a_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l226_c267_c80a_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l226_c237_7f8b_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l226_c207_e041_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l226_c176_f437_return_output, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l297_c43_4a0d_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l296_c17_3517 := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c40_e9c0_return_output.data;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l296_c17_3517;
     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded[chacha20poly1305_decrypt_tb_c_l226_c108_8ded] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_chacha20poly1305_decrypt_tb_c_l226_c108_8ded_arg3;
     -- Outputs

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l280_c9_0d90] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l294_c13_1fd5] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;

     -- Submodule level 8
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_0d90_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l294_c13_1fd5_return_output;
     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l280_c9_1dc0] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l291_c9_3854] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;

     -- Submodule level 9
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l280_c9_1dc0_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l291_c9_3854_return_output;
     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l281_c1_6d2f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l280_c5_af52] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;

     -- Submodule level 10
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l281_c1_6d2f_return_output;
     REG_VAR_ciphertext_in_stream := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     REG_VAR_ciphertext_remaining_in := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     REG_VAR_output_packet_count := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     REG_VAR_plaintext_out_expected := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     REG_VAR_plaintext_out_size := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     REG_VAR_plaintext_remaining_out := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l280_c5_af52_return_output;
     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l313_c9_a764] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l283_c1_dfa4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l292_c1_22cd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l285_c1_5a6d] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output;

     -- Submodule level 11
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l313_c9_a764_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l285_c1_5a6d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l283_c1_dfa4_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l292_c1_22cd_return_output;
     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l313_c5_fec8] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a[chacha20poly1305_decrypt_tb_c_l284_c13_746a] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l284_c13_746a_chacha20poly1305_decrypt_tb_c_l284_c13_746a_arg0;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l294_c1_fccf] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f[chacha20poly1305_decrypt_tb_c_l286_c13_4b4f] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_chacha20poly1305_decrypt_tb_c_l286_c13_4b4f_arg0;
     -- Outputs

     -- Submodule level 12
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l294_c1_fccf_return_output;
     REG_VAR_tag_match_checked := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l313_c5_fec8_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7[chacha20poly1305_decrypt_tb_c_l298_c17_f8d7] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_chacha20poly1305_decrypt_tb_c_l298_c17_f8d7_arg1;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274[chacha20poly1305_decrypt_tb_c_l306_c17_8274] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l306_c17_8274_chacha20poly1305_decrypt_tb_c_l306_c17_8274_arg1;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_input_packet_count <= REG_VAR_input_packet_count;
REG_COMB_ciphertext_in_stream <= REG_VAR_ciphertext_in_stream;
REG_COMB_ciphertext_remaining_in <= REG_VAR_ciphertext_remaining_in;
REG_COMB_cycle_counter <= REG_VAR_cycle_counter;
REG_COMB_output_packet_count <= REG_VAR_output_packet_count;
REG_COMB_plaintext_out_size <= REG_VAR_plaintext_out_size;
REG_COMB_plaintext_remaining_out <= REG_VAR_plaintext_remaining_out;
REG_COMB_plaintext_out_expected <= REG_VAR_plaintext_out_expected;
REG_COMB_tag_match_checked <= REG_VAR_tag_match_checked;
REG_COMB_chacha20poly1305_decrypt_axis_in <= REG_VAR_chacha20poly1305_decrypt_axis_in;
-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_key <= VAR_chacha20poly1305_decrypt_key;
else
  module_to_global.chacha20poly1305_decrypt_key <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_nonce <= VAR_chacha20poly1305_decrypt_nonce;
else
  module_to_global.chacha20poly1305_decrypt_nonce <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad <= VAR_chacha20poly1305_decrypt_aad;
else
  module_to_global.chacha20poly1305_decrypt_aad <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad_len <= VAR_chacha20poly1305_decrypt_aad_len;
else
  module_to_global.chacha20poly1305_decrypt_aad_len <= to_unsigned(0, 8);
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= VAR_chacha20poly1305_decrypt_axis_out_ready;
else
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     input_packet_count <= REG_COMB_input_packet_count;
     ciphertext_in_stream <= REG_COMB_ciphertext_in_stream;
     ciphertext_remaining_in <= REG_COMB_ciphertext_remaining_in;
     cycle_counter <= REG_COMB_cycle_counter;
     output_packet_count <= REG_COMB_output_packet_count;
     plaintext_out_size <= REG_COMB_plaintext_out_size;
     plaintext_remaining_out <= REG_COMB_plaintext_remaining_out;
     plaintext_out_expected <= REG_COMB_plaintext_out_expected;
     tag_match_checked <= REG_COMB_tag_match_checked;
     chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in;
 end if;
 end if;
end process;
-- Shared global regs
module_to_global.chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in when clk_en_internal='1' else chacha20poly1305_decrypt_axis_in;

end arch;
