//==========================================================================
// Copyright (C) 2024 Chili.CHIPS*ba
//--------------------------------------------------------------------------
//                      PROPRIETARY INFORMATION
//
// The information contained in this file is the property of CHILI CHIPS LLC.
// Except as specifically authorized in writing by CHILI CHIPS LLC, the holder
// of this file: (1) shall keep all information contained herein confidential;
// and (2) shall protect the same in whole or in part from disclosure and
// dissemination to all third parties; and (3) shall use the same for operation
// and maintenance purposes only.
//--------------------------------------------------------------------------
// Description: 
//   DPE Multiplexer
//==========================================================================

module dpe_multiplexer #(
    parameter TDATA_WIDTH = 128,
    parameter TUSER_WIDTH = 5
) (
    input  logic      clk,
    input  logic      rst,
    
    input  logic      pause,
    output logic      is_idle,
    
    dpe_if.s_axis     inp0,
    dpe_if.s_axis     inp1,
    dpe_if.s_axis     inp2,
    dpe_if.s_axis     inp3,
    dpe_if.s_axis     inp4,
    dpe_if.m_axis     outp
);
    typedef enum logic [3:0] {
        IDLE,
        R0, S0,
        R1, S1,
        R2, S2,
        R3, S3,
        R4, S4
    } state_t;
    
    state_t state, next_state;
    
    logic                          s_tready;
    logic                          s_tvalid;
    logic [TDATA_WIDTH-1:0]        s_tdata;
    logic                          s_tlast;
    logic [(TDATA_WIDTH+7)/8-1:0]  s_tkeep;
    logic [TUSER_WIDTH-1:0]        s_tuser;
    logic                          s_out_tvalid;
    
    // FSM registers
    always_ff @(posedge clk) begin
        if (rst) begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end
    
    // FSM transition logic
    always_comb begin
        next_state = state;
        
        case (state)
            IDLE: begin
                if (!pause) next_state = R0;
            end
            
            R0: begin
                if (inp0.tvalid && s_tready)         next_state = S0;
                else if (pause)                      next_state = IDLE;
                else if (!inp0.tvalid && s_tready)   next_state = R1;
            end
            
            S0: begin
                if (inp0.tlast && inp0.tvalid && s_tready) begin
                    next_state = pause ? IDLE : R1;
                end
            end
            
            R1: begin
                if (inp1.tvalid && s_tready)         next_state = S1;
                else if (pause)                      next_state = IDLE;
                else if (!inp1.tvalid && s_tready)   next_state = R2;
            end
            
            S1: begin
                if (inp1.tlast && inp1.tvalid && s_tready) begin
                    next_state = pause ? IDLE : R2;
                end
            end
            
            R2: begin
                if (inp2.tvalid && s_tready)         next_state = S2;
                else if (pause)                      next_state = IDLE;
                else if (!inp2.tvalid && s_tready)   next_state = R3;
            end
            
            S2: begin
                if (inp2.tlast && inp2.tvalid && s_tready) begin
                    next_state = pause ? IDLE : R3;
                end
            end
            
            R3: begin
                if (inp3.tvalid && s_tready)         next_state = S3;
                else if (pause)                      next_state = IDLE;
                else if (!inp3.tvalid && s_tready)   next_state = R4;
            end
            
            S3: begin
                if (inp3.tlast && inp3.tvalid && s_tready) begin
                    next_state = pause ? IDLE : R4;
                end
            end
            
            R4: begin
                if (inp4.tvalid && s_tready)         next_state = S4;
                else if (pause)                      next_state = IDLE;
                else if (!inp4.tvalid && s_tready)   next_state = R0;
            end
            
            S4: begin
                if (inp4.tlast && inp4.tvalid && s_tready) begin
                    next_state = pause ? IDLE : R0;
                end
            end
            
            default:
                next_state = state;
        endcase
    end
    
    // Outputs logic
    always_comb begin
        // Default assignments
        is_idle = 0;
        s_tvalid = 0;
        s_tdata = '0;
        s_tlast = 0;
        s_tkeep = '0;
        s_tuser = '0;
        inp0.tready = 0;
        inp1.tready = 0;
        inp2.tready = 0;
        inp3.tready = 0;
        inp4.tready = 0;
        
        case (state)
            IDLE: begin
                is_idle = !s_out_tvalid;
            end
            
            R0, S0: begin
                is_idle = 0;
                s_tvalid = inp0.tvalid;
                s_tdata = inp0.tdata;
                s_tlast = inp0.tlast;
                s_tkeep = inp0.tkeep;
                s_tuser = 5'b00001;
                inp0.tready = s_tready;
            end
            
            R1, S1: begin
                is_idle = 0;
                s_tvalid = inp1.tvalid;
                s_tdata = inp1.tdata;
                s_tlast = inp1.tlast;
                s_tkeep = inp1.tkeep;
                s_tuser = 5'b00010;
                inp1.tready = s_tready;
            end
            
            R2, S2: begin
                is_idle = 0;
                s_tvalid = inp2.tvalid;
                s_tdata = inp2.tdata;
                s_tlast = inp2.tlast;
                s_tkeep = inp2.tkeep;
                s_tuser = 5'b00100;
                inp2.tready = s_tready;
            end
            
            R3, S3: begin
                is_idle = 0;
                s_tvalid = inp3.tvalid;
                s_tdata = inp3.tdata;
                s_tlast = inp3.tlast;
                s_tkeep = inp3.tkeep;
                s_tuser = 5'b01000;
                inp3.tready = s_tready;
            end
            
            R4, S4: begin
                is_idle = 0;
                s_tvalid = inp4.tvalid;
                s_tdata = inp4.tdata;
                s_tlast = inp4.tlast;
                s_tkeep = inp4.tkeep;
                s_tuser = 5'b10000;
                inp4.tready = s_tready;
            end
            
            default:
                is_idle = !s_out_tvalid;
        endcase
    end
    
    assign outp.tvalid = s_out_tvalid;
    
    // Skid buffer
    axis_register #(
        .DATA_WIDTH(TDATA_WIDTH),
        .USER_WIDTH(TUSER_WIDTH)
    ) sbuff (
        .clk(clk),
        .rst(rst),
        .s_axis_tvalid(s_tvalid),
        .s_axis_tready(s_tready),
        .s_axis_tdata(s_tdata),
        .s_axis_tkeep(s_tkeep),
        .s_axis_tlast(s_tlast),
        .s_axis_tuser(s_tuser),
        .s_axis_tid('0),
        .s_axis_tdest('0),
        .m_axis_tvalid(s_out_tvalid),
        .m_axis_tready(outp.tready),
        .m_axis_tdata(outp.tdata),
        .m_axis_tkeep(outp.tkeep),
        .m_axis_tlast(outp.tlast),
        .m_axis_tuser(outp.tuser),
        .m_axis_tid(),
        .m_axis_tdest()
    );
endmodule
