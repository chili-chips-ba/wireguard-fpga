-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.8059474611482419]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_db8fd939 is
port(
 clk : in std_logic;
 elem_val : in unsigned(31 downto 0);
 ref_toks_0 : in chacha20_state;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint32_t_array_16_t);
end VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_db8fd939;
architecture arch of VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_1CLK_db8fd939 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 1;
-- All of the wires/regs in function
-- Stage 0
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse : unsigned(31 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse : unsigned(31 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse : unsigned(31 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse : unsigned(31 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse : unsigned(31 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse : unsigned(31 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse : unsigned(31 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse : unsigned(31 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse : unsigned(31 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse : unsigned(31 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse : unsigned(31 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse : unsigned(31 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse : unsigned(31 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse : unsigned(31 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse : unsigned(31 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse : unsigned(31 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint32_t_array_16_t is
 
  variable base : uint32_t_array_16_t; 
  variable return_output : uint32_t_array_16_t;
begin
      base.data(2) := ref_toks_0;
      base.data(5) := ref_toks_1;
      base.data(11) := ref_toks_2;
      base.data(8) := ref_toks_3;
      base.data(14) := ref_toks_4;
      base.data(0) := ref_toks_5;
      base.data(3) := ref_toks_6;
      base.data(9) := ref_toks_7;
      base.data(6) := ref_toks_8;
      base.data(12) := ref_toks_9;
      base.data(15) := ref_toks_10;
      base.data(4) := ref_toks_11;
      base.data(1) := ref_toks_12;
      base.data(7) := ref_toks_13;
      base.data(10) := ref_toks_14;
      base.data(13) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66 : 1 clocks latency
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_b981834f port map (
clk,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef : 1 clocks latency
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da : 1 clocks latency
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459 : 1 clocks latency
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d : 1 clocks latency
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223 : 1 clocks latency
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_4d6d6521 port map (
clk,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8 : 1 clocks latency
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_b981834f port map (
clk,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7 : 1 clocks latency
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32 : 1 clocks latency
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2 : 1 clocks latency
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a : 1 clocks latency
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436 : 1 clocks latency
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75 : 1 clocks latency
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_4d6d6521 port map (
clk,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79 : 1 clocks latency
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016 : 1 clocks latency
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016 : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5 : 0 clocks latency
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb : 1 clocks latency
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb : entity work.MUX_uint1_t_uint32_t_uint32_t_1CLK_6d084181 port map (
clk,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- Registers
 -- Stage 0
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(31 downto 0);
 variable VAR_ref_toks_0 : chacha20_state;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint32_t_array_16_t;
 variable VAR_base : chacha20_state;
 variable VAR_rv : uint32_t_array_16_t;
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5817_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_d228_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c16_c037_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b2a5_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_9c47_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_fca0_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_916b_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_6aaa_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_1c61_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_0858_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_72a3_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_3f3d_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_4985_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_3905_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c16_f28c_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_201e_return_output : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output : unsigned(31 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_409e_return_output : uint32_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right := to_unsigned(14, 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left := VAR_var_dim_0;
     -- CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_1c61] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_1c61_return_output := VAR_ref_toks_0.state(6);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_4985] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_4985_return_output := VAR_ref_toks_0.state(1);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b2a5] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b2a5_return_output := VAR_ref_toks_0.state(8);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c16_c037] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c16_c037_return_output := VAR_ref_toks_0.state(11);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_3f3d] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_3f3d_return_output := VAR_ref_toks_0.state(4);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_201e] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_201e_return_output := VAR_ref_toks_0.state(13);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_9c47] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_9c47_return_output := VAR_ref_toks_0.state(14);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_6aaa] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_6aaa_return_output := VAR_ref_toks_0.state(9);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_fca0] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_fca0_return_output := VAR_ref_toks_0.state(0);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_d228] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_d228_return_output := VAR_ref_toks_0.state(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_72a3] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_72a3_return_output := VAR_ref_toks_0.state(15);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_3905] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_3905_return_output := VAR_ref_toks_0.state(7);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_916b] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_916b_return_output := VAR_ref_toks_0.state(3);

     -- CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c16_f28c] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c16_f28c_return_output := VAR_ref_toks_0.state(10);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_0858] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_0858_return_output := VAR_ref_toks_0.state(12);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output;

     -- CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5817] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5817_return_output := VAR_ref_toks_0.state(2);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output;

     -- Submodule level 1
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l101_c5_a7d4_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l107_c5_f4e6_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l113_c5_fc18_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l119_c5_5344_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l125_c5_6fa5_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l35_c5_96f4_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l41_c5_9e0f_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l47_c5_18e0_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l53_c5_8973_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l59_c5_c7a3_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l65_c5_95ef_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l71_c5_c880_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l77_c5_1b7e_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l83_c5_2278_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l89_c5_a99a_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l95_c5_7e23_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l22_c15_fca0_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l31_c16_f28c_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l19_c16_c037_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l26_c16_0858_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l32_c16_201e_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l21_c16_9c47_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l27_c16_72a3_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l29_c15_4985_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l17_c15_5817_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l23_c15_916b_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l28_c15_3f3d_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l18_c15_d228_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l25_c15_1c61_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l30_c15_3905_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l20_c15_b2a5_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse := VAR_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l24_c15_6aaa_return_output;
     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7] LATENCY=1
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_iffalse;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79] LATENCY=1
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_iffalse;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436] LATENCY=1
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_iffalse;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d] LATENCY=1
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_iffalse;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66] LATENCY=1
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_iffalse;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32] LATENCY=1
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_iffalse;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75] LATENCY=1
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_iffalse;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da] LATENCY=1
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_iffalse;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459] LATENCY=1
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_iffalse;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2] LATENCY=1
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_iffalse;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8] LATENCY=1
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_iffalse;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016] LATENCY=1
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_iffalse;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb] LATENCY=1
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_iffalse;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a] LATENCY=1
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_iffalse;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef] LATENCY=1
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_iffalse;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223] LATENCY=1
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_iffalse;

     -- Write to comb signals
   elsif STAGE = 1 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb[VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_409e] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_409e_return_output := CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb(
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l34_c2_5a66_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l40_c2_30ef_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l46_c2_54da_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l52_c2_9459_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l58_c2_bf1d_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l64_c2_f223_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l70_c2_06a8_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l76_c2_a8f7_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l82_c2_aa32_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l88_c2_f1e2_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l94_c2_059a_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l100_c2_6436_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l106_c2_cc75_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l112_c2_eb79_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l118_c2_9016_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l124_c2_b6eb_return_output);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_uint32_t_array_16_t_uint32_t_array_16_t_b3fb_VAR_REF_ASSIGN_uint32_t_chacha20_state_state_VAR_23da_c_l131_c10_409e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
 end if;
end process;

end arch;
