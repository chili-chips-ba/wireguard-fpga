-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.023255813953488372, 0.046511627906976744, 0.06976744186046512, 0.09302325581395349, 0.11627906976744186, 0.13953488372093023, 0.16279069767441862, 0.18604651162790697, 0.20930232558139533, 0.2325581395348837, 0.25581395348837205, 0.2790697674418604, 0.30232558139534876, 0.3255813953488371, 0.3488372093023255, 0.37209302325581384, 0.3953488372093022, 0.41860465116279055, 0.4418604651162789, 0.46511627906976727, 0.4883720930232556, 0.511627906976744, 0.5348837209302324, 0.5581395348837208, 0.5813953488372092, 0.6046511627906976, 0.627906976744186, 0.6511627906976745, 0.6744186046511629, 0.6976744186046513, 0.7209302325581397, 0.7441860465116281, 0.7674418604651165, 0.790697674418605, 0.8139534883720934, 0.8372093023255818, 0.8604651162790702, 0.8837209302325586, 0.906976744186047, 0.9302325581395354, 0.9534883720930238, 0.9767441860465123]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 3
entity chacha20_decrypt_pipeline_no_handshake_42CLK_cb4da253 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in chacha20_decrypt_pipeline_no_handshake_global_to_module_t;
 module_to_global : out chacha20_decrypt_pipeline_no_handshake_module_to_global_t);
end chacha20_decrypt_pipeline_no_handshake_42CLK_cb4da253;
architecture arch of chacha20_decrypt_pipeline_no_handshake_42CLK_cb4da253 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 42;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 1
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 2
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 3
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 4
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 5
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 6
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 7
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 8
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 9
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 10
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 11
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 12
signal REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 13
signal REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 14
signal REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 15
signal REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 16
signal REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 17
signal REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 18
signal REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 19
signal REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 20
signal REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 21
signal REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 22
signal REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 23
signal REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 24
signal REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 25
signal REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 26
signal REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 27
signal REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 28
signal REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 29
signal REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 30
signal REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 31
signal REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 32
signal REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 33
signal REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 34
signal REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 35
signal REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 36
signal REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 37
signal REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 38
signal REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 39
signal REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 40
signal REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 41
signal REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- chacha20_decrypt_pipeline_no_handshake_in_reg_func[chacha20_decrypt_c_l24_c102_2533]
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data : chacha20_decrypt_loop_body_in_t;
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id : unsigned(7 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output : chacha20_decrypt_pipeline_no_handshake_in_reg_t;

-- chacha20_decrypt_loop_body[chacha20_decrypt_c_l24_c308_83cc]
signal chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs : chacha20_decrypt_loop_body_in_t;
signal chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output : axis512_t;

-- chacha20_decrypt_pipeline_no_handshake_out_reg_func[chacha20_decrypt_c_l24_c397_29e7]
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data : axis512_t;
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output : chacha20_decrypt_pipeline_no_handshake_out_reg_t;


begin

-- SUBMODULE INSTANCES 
-- chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533 : 0 clocks latency
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533 : entity work.chacha20_decrypt_pipeline_no_handshake_in_reg_func_0CLK_b45f1687 port map (
clk,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output);

-- chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc : 42 clocks latency
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc : entity work.chacha20_decrypt_loop_body_42CLK_addc024f port map (
clk,
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs,
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output);

-- chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7 : 0 clocks latency
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7 : entity work.chacha20_decrypt_pipeline_no_handshake_out_reg_func_0CLK_b45f1687 port map (
clk,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 -- Stage 0
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 1
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 2
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 3
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 4
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 5
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 6
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 7
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 8
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 9
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 10
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 11
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 12
 REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 13
 REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 14
 REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 15
 REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 16
 REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 17
 REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 18
 REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 19
 REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 20
 REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 21
 REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 22
 REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 23
 REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 24
 REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 25
 REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 26
 REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 27
 REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 28
 REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 29
 REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 30
 REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 31
 REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 32
 REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 33
 REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 34
 REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 35
 REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 36
 REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 37
 REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 38
 REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 39
 REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 40
 REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Stage 41
 REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id,
 REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid,
 REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output,
 chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output,
 chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_valid : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out : axis512_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_valid : unsigned(0 downto 0);
 variable VAR_i : chacha20_decrypt_pipeline_no_handshake_in_reg_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output : chacha20_decrypt_pipeline_no_handshake_in_reg_t;
 variable VAR_d : axis512_t;
 variable VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs : chacha20_decrypt_loop_body_in_t;
 variable VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_7a3a_return_output : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output : axis512_t;
 variable VAR_o : chacha20_decrypt_pipeline_no_handshake_out_reg_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data : axis512_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_dbec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_e940_return_output : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output : chacha20_decrypt_pipeline_no_handshake_out_reg_t;
 variable VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_4b77_return_output : axis512_t;
 variable VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_0991_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_64d6_return_output : unsigned(0 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id := to_unsigned(0, 8);
 -- Reads from global variables
     VAR_chacha20_decrypt_pipeline_no_handshake_in := global_to_module.chacha20_decrypt_pipeline_no_handshake_in;
     VAR_chacha20_decrypt_pipeline_no_handshake_in_valid := global_to_module.chacha20_decrypt_pipeline_no_handshake_in_valid;
     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid := VAR_chacha20_decrypt_pipeline_no_handshake_in_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data := VAR_chacha20_decrypt_pipeline_no_handshake_in;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     -- chacha20_decrypt_pipeline_no_handshake_in_reg_func[chacha20_decrypt_c_l24_c102_2533] LATENCY=0
     -- Clock enable
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_CLOCK_ENABLE;
     -- Inputs
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_data;
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_id;
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_valid;
     -- Outputs
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output := chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d[chacha20_decrypt_c_l24_c459_e940] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_e940_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output.valid;

     -- CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d[chacha20_decrypt_c_l24_c453_dbec] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_dbec_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output.id;

     -- CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d[chacha20_decrypt_c_l24_c335_7a3a] LATENCY=0
     VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_7a3a_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_2533_return_output.data;

     -- Submodule level 2
     VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs := VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_7a3a_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_e940_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_dbec_return_output;
     -- chacha20_decrypt_loop_body[chacha20_decrypt_c_l24_c308_83cc] LATENCY=42
     -- Inputs
     chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs <= VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_inputs;

     -- Write to comb signals
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 26 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 27 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 28 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 29 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 30 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 31 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 32 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 33 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 34 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 35 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 36 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 37 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 38 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 39 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 40 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 41 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
   elsif STAGE = 42 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id := REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid := REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE := REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Submodule outputs
     VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output := chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output;

     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data := VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_83cc_return_output;
     -- chacha20_decrypt_pipeline_no_handshake_out_reg_func[chacha20_decrypt_c_l24_c397_29e7] LATENCY=0
     -- Clock enable
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Inputs
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_data;
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     -- Outputs
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output := chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d[chacha20_decrypt_c_l24_c515_4b77] LATENCY=0
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_4b77_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output.data;

     -- CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d[chacha20_decrypt_c_l24_c571_0991] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_0991_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output.id;

     -- CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d[chacha20_decrypt_c_l24_c628_64d6] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_64d6_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_return_output.valid;

     -- Submodule level 2
     VAR_chacha20_decrypt_pipeline_no_handshake_out := VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_4b77_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_valid := VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_64d6_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_id := VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_0991_return_output;
   end if;
 end loop;

-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out <= VAR_chacha20_decrypt_pipeline_no_handshake_out;
else
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out <= axis512_t_NULL;
end if;
if clk_en_internal='1' then
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_valid;
else
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out_valid <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     -- Stage 0
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 1
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 2
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 3
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 4
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 5
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 6
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 7
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 8
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 9
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 10
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 11
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 12
     REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE12_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 13
     REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE13_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 14
     REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE14_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 15
     REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE15_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 16
     REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE16_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 17
     REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE17_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 18
     REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE18_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 19
     REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE19_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 20
     REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE20_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 21
     REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE21_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 22
     REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE22_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 23
     REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE23_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 24
     REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE24_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 25
     REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE25_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 26
     REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE26_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 27
     REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE27_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 28
     REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE28_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 29
     REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE29_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 30
     REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE30_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 31
     REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE31_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 32
     REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE32_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 33
     REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE33_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 34
     REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE34_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 35
     REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE35_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 36
     REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE36_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 37
     REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE37_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 38
     REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE38_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 39
     REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE39_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 40
     REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE40_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
     -- Stage 41
     REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id <= COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_id;
     REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid <= COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_valid;
     REG_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE <= COMB_STAGE41_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_29e7_CLOCK_ENABLE;
 end if;
 end if;
end process;

end arch;
