-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 6
entity u320_t_to_bytes_0CLK_801a240b is
port(
 x : in u320_t;
 return_output : out uint8_t_array_40_t);
end u320_t_to_bytes_0CLK_801a240b;
architecture arch of u320_t_to_bytes_0CLK_801a240b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd]
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd]
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd]
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd]
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd]
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
signal FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;

function CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned) return uint8_t_array_40_t is
 
  variable base : uint8_t_array_40_t; 
  variable return_output : uint8_t_array_40_t;
begin
      base.data(0) := ref_toks_0;
      base.data(1) := ref_toks_1;
      base.data(2) := ref_toks_2;
      base.data(3) := ref_toks_3;
      base.data(4) := ref_toks_4;
      base.data(5) := ref_toks_5;
      base.data(6) := ref_toks_6;
      base.data(7) := ref_toks_7;
      base.data(8) := ref_toks_8;
      base.data(9) := ref_toks_9;
      base.data(10) := ref_toks_10;
      base.data(11) := ref_toks_11;
      base.data(12) := ref_toks_12;
      base.data(13) := ref_toks_13;
      base.data(14) := ref_toks_14;
      base.data(15) := ref_toks_15;
      base.data(16) := ref_toks_16;
      base.data(17) := ref_toks_17;
      base.data(18) := ref_toks_18;
      base.data(19) := ref_toks_19;
      base.data(20) := ref_toks_20;
      base.data(21) := ref_toks_21;
      base.data(22) := ref_toks_22;
      base.data(23) := ref_toks_23;
      base.data(24) := ref_toks_24;
      base.data(25) := ref_toks_25;
      base.data(26) := ref_toks_26;
      base.data(27) := ref_toks_27;
      base.data(28) := ref_toks_28;
      base.data(29) := ref_toks_29;
      base.data(30) := ref_toks_30;
      base.data(31) := ref_toks_31;
      base.data(32) := ref_toks_32;
      base.data(33) := ref_toks_33;
      base.data(34) := ref_toks_34;
      base.data(35) := ref_toks_35;
      base.data(36) := ref_toks_36;
      base.data(37) := ref_toks_37;
      base.data(38) := ref_toks_38;
      base.data(39) := ref_toks_39;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : 0 clocks latency
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : entity work.uint64_t_to_bytes_0CLK_25f4cd11 port map (
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x,
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output);

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : 0 clocks latency
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : entity work.uint64_t_to_bytes_0CLK_25f4cd11 port map (
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x,
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output);

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : 0 clocks latency
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : entity work.uint64_t_to_bytes_0CLK_25f4cd11 port map (
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x,
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output);

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : 0 clocks latency
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : entity work.uint64_t_to_bytes_0CLK_25f4cd11 port map (
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x,
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output);

-- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : 0 clocks latency
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd : entity work.uint64_t_to_bytes_0CLK_25f4cd11 port map (
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x,
FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 x,
 -- All submodule outputs
 FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output,
 FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output,
 FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output,
 FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output,
 FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : uint8_t_array_40_t;
 variable VAR_x : u320_t;
 variable VAR_rv : uint8_t_array_40_t;
 variable VAR_pos : unsigned(6 downto 0);
 variable VAR_field_pos : unsigned(6 downto 0);
 variable VAR_limbs_dim_0 : unsigned(2 downto 0);
 variable VAR_limbs_elem_bytes : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output : unsigned(63 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output : uint8_t_array_8_t;
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb_u320_t_bytes_t_h_l25_c12_1a6e_return_output : uint8_t_array_40_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_x := x;

     -- Submodule level 0
     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[u320_t_bytes_t_h_l17_c57_6000] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output := VAR_x.limbs(3);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[u320_t_bytes_t_h_l17_c57_6000] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output := VAR_x.limbs(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[u320_t_bytes_t_h_l17_c57_6000] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output := VAR_x.limbs(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[u320_t_bytes_t_h_l17_c57_6000] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output := VAR_x.limbs(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[u320_t_bytes_t_h_l17_c57_6000] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output := VAR_x.limbs(4);

     -- Submodule level 1
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output;
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output;
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output;
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output;
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_u320_t_bytes_t_h_l17_c57_6000_return_output;
     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x <= VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output := FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output;

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x <= VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output := FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output;

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x <= VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output := FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output;

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x <= VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output := FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output;

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes[u320_t_bytes_t_h_l17_c39_accd] LATENCY=0
     -- Inputs
     FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x <= VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_x;
     -- Outputs
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output := FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output;

     -- Submodule level 2
     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(4);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(4);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(3);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(7);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(5);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(5);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(4);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(5);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(4);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(5);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(6);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(6);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(5);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(6);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(2);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(6);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(7);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(3);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(3);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(4);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(7);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(7);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(3);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(7);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(6);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(0);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(1);

     -- FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d[u320_t_bytes_t_h_l20_c20_8cbc] LATENCY=0
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output := VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_uint64_t_to_bytes_u320_t_bytes_t_h_l17_c39_accd_return_output.data(3);

     -- Submodule level 3
     -- CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb[u320_t_bytes_t_h_l25_c12_1a6e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb_u320_t_bytes_t_h_l25_c12_1a6e_return_output := CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb(
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_0_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_1_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_2_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_3_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_0_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_1_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_2_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_3_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_4_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_4_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_5_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_5_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_6_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_6_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output,
     VAR_FOR_u320_t_bytes_t_h_l16_c1_184d_ITER_4_FOR_u320_t_bytes_t_h_l18_c2_0fbe_ITER_7_CONST_REF_RD_uint8_t_uint8_t_array_8_t_data_7_d41d_u320_t_bytes_t_h_l20_c20_8cbc_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_40_t_uint8_t_array_40_t_54cb_u320_t_bytes_t_h_l25_c12_1a6e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
