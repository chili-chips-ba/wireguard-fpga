-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.20810055865921787, 0.5921787709497207, 0.9762569832402235]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_3CLK_087b5579 is
port(
 clk : in std_logic;
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_3CLK_087b5579;
architecture arch of uint320_mul_3CLK_087b5579 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 3;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
-- Stage 1
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
-- Stage 2
signal REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_7657]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_93c2]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_ae83]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_2807]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_8adc]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_07e1]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_39b7]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_979f]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_6054]
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d81e]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8f19]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6117]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_8fbd]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_5ab2]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_f2b2]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_7183]
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_ecf7]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_1680]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6982]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_395c]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_b94d]
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_f995]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_eeeb]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_4363]
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15]
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c]
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_3b5f]
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_9ca18c4f port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_eec62983 port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right,
FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd : entity work.BIN_OP_PLUS_uint64_t_uint1_t_1CLK_9324e8e6 port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0f464748 port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right,
FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_ec635a74 port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7 : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0320092f port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right,
FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right,
FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : 0 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output);

-- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f : 1 clocks latency
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_8f2211ba port map (
clk,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right,
FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- Registers
 -- Stage 0
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 -- Stage 1
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left,
 -- Stage 2
 REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output,
 FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_ccca_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_ccca_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_ccca_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_ccca_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_a867_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_ccca_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_e5a8_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_73b7_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_a867_DUPLICATE_2e26_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_a867_DUPLICATE_4110_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_e301_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_645d_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse := to_unsigned(0, 64);
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_ccca] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_ccca_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_ccca] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_ccca_return_output := u320_t_NULL.limbs(1);

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_ccca] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_ccca_return_output := u320_t_NULL.limbs(2);

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_ccca] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_ccca_return_output := u320_t_NULL.limbs(0);

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_ccca] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_ccca_return_output := u320_t_NULL.limbs(4);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_ccca_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_ccca_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_ccca_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_ccca_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_ccca_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_e5a8]_DUPLICATE_645d LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_645d_return_output := VAR_a.limbs(3);

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_a867] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_a867_return_output := VAR_b.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_e5a8]_DUPLICATE_e301 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_e301_return_output := VAR_a.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_a867]_DUPLICATE_17b8 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output := VAR_b.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_a867]_DUPLICATE_4110 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_a867_DUPLICATE_4110_return_output := VAR_b.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_a867]_DUPLICATE_1c3b LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_a867]_DUPLICATE_2e26 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_a867_DUPLICATE_2e26_return_output := VAR_b.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_e5a8]_DUPLICATE_bb80 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output := VAR_a.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_e5a8]_DUPLICATE_2bc0 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output := VAR_a.limbs(1);

     -- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_e5a8] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_e5a8_return_output := VAR_a.limbs(4);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_bb80_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_a867_DUPLICATE_17b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_2bc0_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_a867_DUPLICATE_1c3b_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_e301_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_e301_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_e301_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_a867_DUPLICATE_2e26_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_a867_DUPLICATE_2e26_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_a867_DUPLICATE_2e26_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_645d_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_e5a8_DUPLICATE_645d_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_a867_DUPLICATE_4110_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_a867_DUPLICATE_4110_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_a867_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_e5a8_return_output;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_2a15] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_2a15_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_product_poly1305_h_l127_c22_6d14_0;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_product_poly1305_h_l127_c22_6d14_0;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_7657] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;

     -- Write to comb signals
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_7657_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l132_c21_1ea9_return_output;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_93c2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_93c2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_ae83] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d81e] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d81e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_2807] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_2807_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_8adc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8f19] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8f19_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6117] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6117_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_07e1] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_07e1_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_39b7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_ecf7] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_8fbd] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_right;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_right;

     -- Write to comb signals
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8fbd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_ecf7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_5ab2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_5ab2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_979f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_6054] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output := FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_1680] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_1680_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_f2b2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6982] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_f2b2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6982_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_7183] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_left;
     FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output := FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_7183_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_f995] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_78d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_f995_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l131_c13_506d;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_b250] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l132_c21_1ea9] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_395c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_395c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_b250_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l132_c21_1ea9_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_high_poly1305_h_l134_c13_38a1;
     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX[poly1305_h_l134_c22_bb97] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_cond;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iftrue;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_b94d] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_left;
     FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output := FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b94d_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_MUX_poly1305_h_l134_c22_bb97_return_output;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_eeeb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eeeb_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_high_poly1305_h_l134_c13_38a1;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_4363] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_left;
     FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output := FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_4363_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right := VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_low_poly1305_h_l133_c13_2064;
     -- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_e96c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output := FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left := VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l131_c13_506d;
     -- FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_3b5f] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_left;
     FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_right;

     -- Write to comb signals
     COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output := FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 := resize(VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_3b5f_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_73b7] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_73b7_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064,
     VAR_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_73b7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_ae83_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_8adc_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_39b7_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     -- Stage 1
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_979f_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_6054_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_78d3_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_c881_ITER_4_FOR_poly1305_h_l123_c9_f216_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_e96c_left;
     -- Stage 2
     REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_0_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_1_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_2_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
     REG_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_c881_ITER_3_FOR_poly1305_h_l123_c9_f216_ITER_0_low_poly1305_h_l133_c13_2064;
 end if;
end process;

end arch;
