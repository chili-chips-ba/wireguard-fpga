
module progmem (
    // Clock & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata,
	// Rewrite firmware
    input  wire        wen,
	input  wire [31:0] waddr,
	input  wire [31:0] wdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 13;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin
    mem['h0000] <= 32'h00000093;
    mem['h0001] <= 32'h00000193;
    mem['h0002] <= 32'h00000213;
    mem['h0003] <= 32'h00000293;
    mem['h0004] <= 32'h00000313;
    mem['h0005] <= 32'h00000393;
    mem['h0006] <= 32'h00000413;
    mem['h0007] <= 32'h00000493;
    mem['h0008] <= 32'h00000513;
    mem['h0009] <= 32'h00000593;
    mem['h000A] <= 32'h00000613;
    mem['h000B] <= 32'h00000693;
    mem['h000C] <= 32'h00000713;
    mem['h000D] <= 32'h00000793;
    mem['h000E] <= 32'h00000813;
    mem['h000F] <= 32'h00000893;
    mem['h0010] <= 32'h00000913;
    mem['h0011] <= 32'h00000993;
    mem['h0012] <= 32'h00000A13;
    mem['h0013] <= 32'h00000A93;
    mem['h0014] <= 32'h00000B13;
    mem['h0015] <= 32'h00000B93;
    mem['h0016] <= 32'h00000C13;
    mem['h0017] <= 32'h00000C93;
    mem['h0018] <= 32'h00000D13;
    mem['h0019] <= 32'h00000D93;
    mem['h001A] <= 32'h00000E13;
    mem['h001B] <= 32'h00000E93;
    mem['h001C] <= 32'h00000F13;
    mem['h001D] <= 32'h00000F93;
    mem['h001E] <= 32'h00000513;
    mem['h001F] <= 32'h00000593;
    mem['h0020] <= 32'h00B52023;
    mem['h0021] <= 32'h00450513;
    mem['h0022] <= 32'hFE254CE3;
    mem['h0023] <= 32'h00001517;
    mem['h0024] <= 32'h3CC50513;
    mem['h0025] <= 32'h00000593;
    mem['h0026] <= 32'h00000613;
    mem['h0027] <= 32'h00C5DC63;
    mem['h0028] <= 32'h00052683;
    mem['h0029] <= 32'h00D5A023;
    mem['h002A] <= 32'h00450513;
    mem['h002B] <= 32'h00458593;
    mem['h002C] <= 32'hFEC5C8E3;
    mem['h002D] <= 32'h00000513;
    mem['h002E] <= 32'h00000593;
    mem['h002F] <= 32'h00B55863;
    mem['h0030] <= 32'h00052023;
    mem['h0031] <= 32'h00450513;
    mem['h0032] <= 32'hFEB54CE3;
    mem['h0033] <= 32'h008000EF;
    mem['h0034] <= 32'h0000006F;
    mem['h0035] <= 32'hFC010113;
    mem['h0036] <= 32'h02112E23;
    mem['h0037] <= 32'h02812C23;
    mem['h0038] <= 32'h04010413;
    mem['h0039] <= 32'hFCC40793;
    mem['h003A] <= 32'h00078513;
    mem['h003B] <= 32'h0A4000EF;
    mem['h003C] <= 32'h06400593;
    mem['h003D] <= 32'h00A00513;
    mem['h003E] <= 32'h1E0000EF;
    mem['h003F] <= 32'hFEA42623;
    mem['h0040] <= 32'h00000793;
    mem['h0041] <= 32'h00078513;
    mem['h0042] <= 32'h03C12083;
    mem['h0043] <= 32'h03812403;
    mem['h0044] <= 32'h04010113;
    mem['h0045] <= 32'h00008067;
    mem['h0046] <= 32'hFE010113;
    mem['h0047] <= 32'h00812E23;
    mem['h0048] <= 32'h02010413;
    mem['h0049] <= 32'hC00027F3;
    mem['h004A] <= 32'hFEF42623;
    mem['h004B] <= 32'hFEC42783;
    mem['h004C] <= 32'h00078513;
    mem['h004D] <= 32'h01C12403;
    mem['h004E] <= 32'h02010113;
    mem['h004F] <= 32'h00008067;
    mem['h0050] <= 32'hFE010113;
    mem['h0051] <= 32'h00812E23;
    mem['h0052] <= 32'h02010413;
    mem['h0053] <= 32'hFE0407A3;
    mem['h0054] <= 32'h01C0006F;
    mem['h0055] <= 32'h00000013;
    mem['h0056] <= 32'hFEF44783;
    mem['h0057] <= 32'h0FF7F793;
    mem['h0058] <= 32'h00178793;
    mem['h0059] <= 32'h0FF7F793;
    mem['h005A] <= 32'hFEF407A3;
    mem['h005B] <= 32'hFEF44783;
    mem['h005C] <= 32'h0FF7F713;
    mem['h005D] <= 32'h00700793;
    mem['h005E] <= 32'hFCE7FEE3;
    mem['h005F] <= 32'h00000013;
    mem['h0060] <= 32'h00000013;
    mem['h0061] <= 32'h01C12403;
    mem['h0062] <= 32'h02010113;
    mem['h0063] <= 32'h00008067;
    mem['h0064] <= 32'hF5010113;
    mem['h0065] <= 32'h0A112623;
    mem['h0066] <= 32'h0A812423;
    mem['h0067] <= 32'h0B010413;
    mem['h0068] <= 32'hF4A42E23;
    mem['h0069] <= 32'hFE042623;
    mem['h006A] <= 32'h0900006F;
    mem['h006B] <= 32'hF6DFF0EF;
    mem['h006C] <= 32'hFEA42423;
    mem['h006D] <= 32'hFE842783;
    mem['h006E] <= 32'h0077D793;
    mem['h006F] <= 32'hFE842703;
    mem['h0070] <= 32'h00F747B3;
    mem['h0071] <= 32'hFEF42423;
    mem['h0072] <= 32'hFE842703;
    mem['h0073] <= 32'h6C0797B7;
    mem['h0074] <= 32'h96578793;
    mem['h0075] <= 32'h02F707B3;
    mem['h0076] <= 32'hFEF42423;
    mem['h0077] <= 32'hFE842783;
    mem['h0078] <= 32'h00B7D793;
    mem['h0079] <= 32'hFE842703;
    mem['h007A] <= 32'h00F747B3;
    mem['h007B] <= 32'hFEF42423;
    mem['h007C] <= 32'hFEC42703;
    mem['h007D] <= 32'h5D5897B7;
    mem['h007E] <= 32'hB6578793;
    mem['h007F] <= 32'h02F707B3;
    mem['h0080] <= 32'h00078713;
    mem['h0081] <= 32'hFE842783;
    mem['h0082] <= 32'h00E787B3;
    mem['h0083] <= 32'hFEF42423;
    mem['h0084] <= 32'hFEC42783;
    mem['h0085] <= 32'h00279793;
    mem['h0086] <= 32'hFF078793;
    mem['h0087] <= 32'h008787B3;
    mem['h0088] <= 32'hFE842703;
    mem['h0089] <= 32'hFAE7AC23;
    mem['h008A] <= 32'hF19FF0EF;
    mem['h008B] <= 32'hFEC42783;
    mem['h008C] <= 32'h00178793;
    mem['h008D] <= 32'hFEF42623;
    mem['h008E] <= 32'hFEC42703;
    mem['h008F] <= 32'h00F00793;
    mem['h0090] <= 32'hF6E7D6E3;
    mem['h0091] <= 32'hFA440793;
    mem['h0092] <= 32'hFAF42223;
    mem['h0093] <= 32'hFA840713;
    mem['h0094] <= 32'hF6040793;
    mem['h0095] <= 32'h04000613;
    mem['h0096] <= 32'h00070593;
    mem['h0097] <= 32'h00078513;
    mem['h0098] <= 32'h7C5000EF;
    mem['h0099] <= 32'hF6040793;
    mem['h009A] <= 32'h04078793;
    mem['h009B] <= 32'hFA440713;
    mem['h009C] <= 32'h00400613;
    mem['h009D] <= 32'h00070593;
    mem['h009E] <= 32'h00078513;
    mem['h009F] <= 32'h7A9000EF;
    mem['h00A0] <= 32'hF6040613;
    mem['h00A1] <= 32'h00000793;
    mem['h00A2] <= 32'h00000713;
    mem['h00A3] <= 32'h04400693;
    mem['h00A4] <= 32'h02000593;
    mem['h00A5] <= 32'hF5C42503;
    mem['h00A6] <= 32'h691000EF;
    mem['h00A7] <= 32'hFA840793;
    mem['h00A8] <= 32'h04000613;
    mem['h00A9] <= 32'h00000593;
    mem['h00AA] <= 32'h00078513;
    mem['h00AB] <= 32'h709000EF;
    mem['h00AC] <= 32'hF6040793;
    mem['h00AD] <= 32'h04400613;
    mem['h00AE] <= 32'h00000593;
    mem['h00AF] <= 32'h00078513;
    mem['h00B0] <= 32'h6F5000EF;
    mem['h00B1] <= 32'h00000013;
    mem['h00B2] <= 32'h0AC12083;
    mem['h00B3] <= 32'h0A812403;
    mem['h00B4] <= 32'h0B010113;
    mem['h00B5] <= 32'h00008067;
    mem['h00B6] <= 32'hFB010113;
    mem['h00B7] <= 32'h04112623;
    mem['h00B8] <= 32'h04812423;
    mem['h00B9] <= 32'h05010413;
    mem['h00BA] <= 32'hFAA42E23;
    mem['h00BB] <= 32'hFAB42C23;
    mem['h00BC] <= 32'hFB842703;
    mem['h00BD] <= 32'hFBC42783;
    mem['h00BE] <= 32'h00E7E663;
    mem['h00BF] <= 32'hFBC42783;
    mem['h00C0] <= 32'h05C0006F;
    mem['h00C1] <= 32'hFD040793;
    mem['h00C2] <= 32'h00078513;
    mem['h00C3] <= 32'hE85FF0EF;
    mem['h00C4] <= 32'hFD040713;
    mem['h00C5] <= 32'hFCC40793;
    mem['h00C6] <= 32'h00400613;
    mem['h00C7] <= 32'h00070593;
    mem['h00C8] <= 32'h00078513;
    mem['h00C9] <= 32'h701000EF;
    mem['h00CA] <= 32'hFD040793;
    mem['h00CB] <= 32'h02000613;
    mem['h00CC] <= 32'h00000593;
    mem['h00CD] <= 32'h00078513;
    mem['h00CE] <= 32'h67D000EF;
    mem['h00CF] <= 32'hFCC42703;
    mem['h00D0] <= 32'hFB842683;
    mem['h00D1] <= 32'hFBC42783;
    mem['h00D2] <= 32'h40F687B3;
    mem['h00D3] <= 32'h00178793;
    mem['h00D4] <= 32'h02F77733;
    mem['h00D5] <= 32'hFBC42783;
    mem['h00D6] <= 32'h00F707B3;
    mem['h00D7] <= 32'h00078513;
    mem['h00D8] <= 32'h04C12083;
    mem['h00D9] <= 32'h04812403;
    mem['h00DA] <= 32'h05010113;
    mem['h00DB] <= 32'h00008067;
    mem['h00DC] <= 32'hEB010113;
    mem['h00DD] <= 32'h14112623;
    mem['h00DE] <= 32'h14812423;
    mem['h00DF] <= 32'h15010413;
    mem['h00E0] <= 32'hEAA42E23;
    mem['h00E1] <= 32'hEAB42C23;
    mem['h00E2] <= 32'h001017B7;
    mem['h00E3] <= 32'h3B878713;
    mem['h00E4] <= 32'hF4C40793;
    mem['h00E5] <= 32'h00070693;
    mem['h00E6] <= 32'h0A000713;
    mem['h00E7] <= 32'h00070613;
    mem['h00E8] <= 32'h00068593;
    mem['h00E9] <= 32'h00078513;
    mem['h00EA] <= 32'h67D000EF;
    mem['h00EB] <= 32'hFE042623;
    mem['h00EC] <= 32'h06C0006F;
    mem['h00ED] <= 32'hEBC42703;
    mem['h00EE] <= 32'hFEC42783;
    mem['h00EF] <= 32'h01078793;
    mem['h00F0] <= 32'h00279793;
    mem['h00F1] <= 32'h00F707B3;
    mem['h00F2] <= 32'h0007A703;
    mem['h00F3] <= 32'hFEC42783;
    mem['h00F4] <= 32'h00279793;
    mem['h00F5] <= 32'hFF078793;
    mem['h00F6] <= 32'h008787B3;
    mem['h00F7] <= 32'hF0E7AE23;
    mem['h00F8] <= 32'hFEC42783;
    mem['h00F9] <= 32'h00878793;
    mem['h00FA] <= 32'h00101737;
    mem['h00FB] <= 32'h39870693;
    mem['h00FC] <= 32'hFEC42703;
    mem['h00FD] <= 32'h00271713;
    mem['h00FE] <= 32'h00E68733;
    mem['h00FF] <= 32'h00072703;
    mem['h0100] <= 32'h00279793;
    mem['h0101] <= 32'hFF078793;
    mem['h0102] <= 32'h008787B3;
    mem['h0103] <= 32'hF0E7AE23;
    mem['h0104] <= 32'hFEC42783;
    mem['h0105] <= 32'h00178793;
    mem['h0106] <= 32'hFEF42623;
    mem['h0107] <= 32'hFEC42703;
    mem['h0108] <= 32'h00700793;
    mem['h0109] <= 32'hF8E7D8E3;
    mem['h010A] <= 32'hF3C42703;
    mem['h010B] <= 32'hEBC42783;
    mem['h010C] <= 32'h0607A783;
    mem['h010D] <= 32'h00F747B3;
    mem['h010E] <= 32'hF2F42E23;
    mem['h010F] <= 32'hF4042703;
    mem['h0110] <= 32'hEBC42783;
    mem['h0111] <= 32'h0647A783;
    mem['h0112] <= 32'h00F747B3;
    mem['h0113] <= 32'hF4F42023;
    mem['h0114] <= 32'hEB842783;
    mem['h0115] <= 32'h00078863;
    mem['h0116] <= 32'hF4442783;
    mem['h0117] <= 32'hFFF7C793;
    mem['h0118] <= 32'hF4F42223;
    mem['h0119] <= 32'hFE042623;
    mem['h011A] <= 32'h09C0006F;
    mem['h011B] <= 32'hFEC42783;
    mem['h011C] <= 32'h00279793;
    mem['h011D] <= 32'hEBC42703;
    mem['h011E] <= 32'h00F707B3;
    mem['h011F] <= 32'h0007C783;
    mem['h0120] <= 32'h00078693;
    mem['h0121] <= 32'hFEC42783;
    mem['h0122] <= 32'h00279793;
    mem['h0123] <= 32'hEBC42703;
    mem['h0124] <= 32'h00F707B3;
    mem['h0125] <= 32'h00178793;
    mem['h0126] <= 32'h0007C783;
    mem['h0127] <= 32'h00879793;
    mem['h0128] <= 32'h00F6C733;
    mem['h0129] <= 32'hFEC42783;
    mem['h012A] <= 32'h00279793;
    mem['h012B] <= 32'hEBC42683;
    mem['h012C] <= 32'h00F687B3;
    mem['h012D] <= 32'h00278793;
    mem['h012E] <= 32'h0007C783;
    mem['h012F] <= 32'h01079793;
    mem['h0130] <= 32'h00F74733;
    mem['h0131] <= 32'hFEC42783;
    mem['h0132] <= 32'h00279793;
    mem['h0133] <= 32'hEBC42683;
    mem['h0134] <= 32'h00F687B3;
    mem['h0135] <= 32'h00378793;
    mem['h0136] <= 32'h0007C783;
    mem['h0137] <= 32'h01879793;
    mem['h0138] <= 32'h00F74733;
    mem['h0139] <= 32'hFEC42783;
    mem['h013A] <= 32'h00279793;
    mem['h013B] <= 32'hFF078793;
    mem['h013C] <= 32'h008787B3;
    mem['h013D] <= 32'hECE7AE23;
    mem['h013E] <= 32'hFEC42783;
    mem['h013F] <= 32'h00178793;
    mem['h0140] <= 32'hFEF42623;
    mem['h0141] <= 32'hFEC42703;
    mem['h0142] <= 32'h00F00793;
    mem['h0143] <= 32'hF6E7D0E3;
    mem['h0144] <= 32'hFE042623;
    mem['h0145] <= 32'h0110006F;
    mem['h0146] <= 32'hF0C42703;
    mem['h0147] <= 32'hF1C42783;
    mem['h0148] <= 32'h00F70733;
    mem['h0149] <= 32'hFEC42783;
    mem['h014A] <= 32'h00479793;
    mem['h014B] <= 32'hFF078793;
    mem['h014C] <= 32'h008787B3;
    mem['h014D] <= 32'hF5C7C783;
    mem['h014E] <= 32'h00279793;
    mem['h014F] <= 32'hFF078793;
    mem['h0150] <= 32'h008787B3;
    mem['h0151] <= 32'hEDC7A783;
    mem['h0152] <= 32'h00F707B3;
    mem['h0153] <= 32'hF0F42623;
    mem['h0154] <= 32'hF3C42703;
    mem['h0155] <= 32'hF0C42783;
    mem['h0156] <= 32'h00F747B3;
    mem['h0157] <= 32'h01079713;
    mem['h0158] <= 32'h0107D793;
    mem['h0159] <= 32'h00E7E7B3;
    mem['h015A] <= 32'hF2F42E23;
    mem['h015B] <= 32'hF2C42703;
    mem['h015C] <= 32'hF3C42783;
    mem['h015D] <= 32'h00F707B3;
    mem['h015E] <= 32'hF2F42623;
    mem['h015F] <= 32'hF1C42703;
    mem['h0160] <= 32'hF2C42783;
    mem['h0161] <= 32'h00F747B3;
    mem['h0162] <= 32'h00C7D713;
    mem['h0163] <= 32'h01479793;
    mem['h0164] <= 32'h00E7E7B3;
    mem['h0165] <= 32'hF0F42E23;
    mem['h0166] <= 32'hF0C42703;
    mem['h0167] <= 32'hF1C42783;
    mem['h0168] <= 32'h00F70733;
    mem['h0169] <= 32'hFEC42783;
    mem['h016A] <= 32'h00479793;
    mem['h016B] <= 32'hFF078793;
    mem['h016C] <= 32'h008787B3;
    mem['h016D] <= 32'hF5D7C783;
    mem['h016E] <= 32'h00279793;
    mem['h016F] <= 32'hFF078793;
    mem['h0170] <= 32'h008787B3;
    mem['h0171] <= 32'hEDC7A783;
    mem['h0172] <= 32'h00F707B3;
    mem['h0173] <= 32'hF0F42623;
    mem['h0174] <= 32'hF3C42703;
    mem['h0175] <= 32'hF0C42783;
    mem['h0176] <= 32'h00F747B3;
    mem['h0177] <= 32'h0087D713;
    mem['h0178] <= 32'h01879793;
    mem['h0179] <= 32'h00E7E7B3;
    mem['h017A] <= 32'hF2F42E23;
    mem['h017B] <= 32'hF2C42703;
    mem['h017C] <= 32'hF3C42783;
    mem['h017D] <= 32'h00F707B3;
    mem['h017E] <= 32'hF2F42623;
    mem['h017F] <= 32'hF1C42703;
    mem['h0180] <= 32'hF2C42783;
    mem['h0181] <= 32'h00F747B3;
    mem['h0182] <= 32'h0077D713;
    mem['h0183] <= 32'h01979793;
    mem['h0184] <= 32'h00E7E7B3;
    mem['h0185] <= 32'hF0F42E23;
    mem['h0186] <= 32'hF1042703;
    mem['h0187] <= 32'hF2042783;
    mem['h0188] <= 32'h00F70733;
    mem['h0189] <= 32'hFEC42783;
    mem['h018A] <= 32'h00479793;
    mem['h018B] <= 32'hFF078793;
    mem['h018C] <= 32'h008787B3;
    mem['h018D] <= 32'hF5E7C783;
    mem['h018E] <= 32'h00279793;
    mem['h018F] <= 32'hFF078793;
    mem['h0190] <= 32'h008787B3;
    mem['h0191] <= 32'hEDC7A783;
    mem['h0192] <= 32'h00F707B3;
    mem['h0193] <= 32'hF0F42823;
    mem['h0194] <= 32'hF4042703;
    mem['h0195] <= 32'hF1042783;
    mem['h0196] <= 32'h00F747B3;
    mem['h0197] <= 32'h01079713;
    mem['h0198] <= 32'h0107D793;
    mem['h0199] <= 32'h00E7E7B3;
    mem['h019A] <= 32'hF4F42023;
    mem['h019B] <= 32'hF3042703;
    mem['h019C] <= 32'hF4042783;
    mem['h019D] <= 32'h00F707B3;
    mem['h019E] <= 32'hF2F42823;
    mem['h019F] <= 32'hF2042703;
    mem['h01A0] <= 32'hF3042783;
    mem['h01A1] <= 32'h00F747B3;
    mem['h01A2] <= 32'h00C7D713;
    mem['h01A3] <= 32'h01479793;
    mem['h01A4] <= 32'h00E7E7B3;
    mem['h01A5] <= 32'hF2F42023;
    mem['h01A6] <= 32'hF1042703;
    mem['h01A7] <= 32'hF2042783;
    mem['h01A8] <= 32'h00F70733;
    mem['h01A9] <= 32'hFEC42783;
    mem['h01AA] <= 32'h00479793;
    mem['h01AB] <= 32'hFF078793;
    mem['h01AC] <= 32'h008787B3;
    mem['h01AD] <= 32'hF5F7C783;
    mem['h01AE] <= 32'h00279793;
    mem['h01AF] <= 32'hFF078793;
    mem['h01B0] <= 32'h008787B3;
    mem['h01B1] <= 32'hEDC7A783;
    mem['h01B2] <= 32'h00F707B3;
    mem['h01B3] <= 32'hF0F42823;
    mem['h01B4] <= 32'hF4042703;
    mem['h01B5] <= 32'hF1042783;
    mem['h01B6] <= 32'h00F747B3;
    mem['h01B7] <= 32'h0087D713;
    mem['h01B8] <= 32'h01879793;
    mem['h01B9] <= 32'h00E7E7B3;
    mem['h01BA] <= 32'hF4F42023;
    mem['h01BB] <= 32'hF3042703;
    mem['h01BC] <= 32'hF4042783;
    mem['h01BD] <= 32'h00F707B3;
    mem['h01BE] <= 32'hF2F42823;
    mem['h01BF] <= 32'hF2042703;
    mem['h01C0] <= 32'hF3042783;
    mem['h01C1] <= 32'h00F747B3;
    mem['h01C2] <= 32'h0077D713;
    mem['h01C3] <= 32'h01979793;
    mem['h01C4] <= 32'h00E7E7B3;
    mem['h01C5] <= 32'hF2F42023;
    mem['h01C6] <= 32'hF1442703;
    mem['h01C7] <= 32'hF2442783;
    mem['h01C8] <= 32'h00F70733;
    mem['h01C9] <= 32'hFEC42783;
    mem['h01CA] <= 32'h00479793;
    mem['h01CB] <= 32'hFF078793;
    mem['h01CC] <= 32'h008787B3;
    mem['h01CD] <= 32'hF607C783;
    mem['h01CE] <= 32'h00279793;
    mem['h01CF] <= 32'hFF078793;
    mem['h01D0] <= 32'h008787B3;
    mem['h01D1] <= 32'hEDC7A783;
    mem['h01D2] <= 32'h00F707B3;
    mem['h01D3] <= 32'hF0F42A23;
    mem['h01D4] <= 32'hF4442703;
    mem['h01D5] <= 32'hF1442783;
    mem['h01D6] <= 32'h00F747B3;
    mem['h01D7] <= 32'h01079713;
    mem['h01D8] <= 32'h0107D793;
    mem['h01D9] <= 32'h00E7E7B3;
    mem['h01DA] <= 32'hF4F42223;
    mem['h01DB] <= 32'hF3442703;
    mem['h01DC] <= 32'hF4442783;
    mem['h01DD] <= 32'h00F707B3;
    mem['h01DE] <= 32'hF2F42A23;
    mem['h01DF] <= 32'hF2442703;
    mem['h01E0] <= 32'hF3442783;
    mem['h01E1] <= 32'h00F747B3;
    mem['h01E2] <= 32'h00C7D713;
    mem['h01E3] <= 32'h01479793;
    mem['h01E4] <= 32'h00E7E7B3;
    mem['h01E5] <= 32'hF2F42223;
    mem['h01E6] <= 32'hF1442703;
    mem['h01E7] <= 32'hF2442783;
    mem['h01E8] <= 32'h00F70733;
    mem['h01E9] <= 32'hFEC42783;
    mem['h01EA] <= 32'h00479793;
    mem['h01EB] <= 32'hFF078793;
    mem['h01EC] <= 32'h008787B3;
    mem['h01ED] <= 32'hF617C783;
    mem['h01EE] <= 32'h00279793;
    mem['h01EF] <= 32'hFF078793;
    mem['h01F0] <= 32'h008787B3;
    mem['h01F1] <= 32'hEDC7A783;
    mem['h01F2] <= 32'h00F707B3;
    mem['h01F3] <= 32'hF0F42A23;
    mem['h01F4] <= 32'hF4442703;
    mem['h01F5] <= 32'hF1442783;
    mem['h01F6] <= 32'h00F747B3;
    mem['h01F7] <= 32'h0087D713;
    mem['h01F8] <= 32'h01879793;
    mem['h01F9] <= 32'h00E7E7B3;
    mem['h01FA] <= 32'hF4F42223;
    mem['h01FB] <= 32'hF3442703;
    mem['h01FC] <= 32'hF4442783;
    mem['h01FD] <= 32'h00F707B3;
    mem['h01FE] <= 32'hF2F42A23;
    mem['h01FF] <= 32'hF2442703;
    mem['h0200] <= 32'hF3442783;
    mem['h0201] <= 32'h00F747B3;
    mem['h0202] <= 32'h0077D713;
    mem['h0203] <= 32'h01979793;
    mem['h0204] <= 32'h00E7E7B3;
    mem['h0205] <= 32'hF2F42223;
    mem['h0206] <= 32'hF1842703;
    mem['h0207] <= 32'hF2842783;
    mem['h0208] <= 32'h00F70733;
    mem['h0209] <= 32'hFEC42783;
    mem['h020A] <= 32'h00479793;
    mem['h020B] <= 32'hFF078793;
    mem['h020C] <= 32'h008787B3;
    mem['h020D] <= 32'hF627C783;
    mem['h020E] <= 32'h00279793;
    mem['h020F] <= 32'hFF078793;
    mem['h0210] <= 32'h008787B3;
    mem['h0211] <= 32'hEDC7A783;
    mem['h0212] <= 32'h00F707B3;
    mem['h0213] <= 32'hF0F42C23;
    mem['h0214] <= 32'hF4842703;
    mem['h0215] <= 32'hF1842783;
    mem['h0216] <= 32'h00F747B3;
    mem['h0217] <= 32'h01079713;
    mem['h0218] <= 32'h0107D793;
    mem['h0219] <= 32'h00E7E7B3;
    mem['h021A] <= 32'hF4F42423;
    mem['h021B] <= 32'hF3842703;
    mem['h021C] <= 32'hF4842783;
    mem['h021D] <= 32'h00F707B3;
    mem['h021E] <= 32'hF2F42C23;
    mem['h021F] <= 32'hF2842703;
    mem['h0220] <= 32'hF3842783;
    mem['h0221] <= 32'h00F747B3;
    mem['h0222] <= 32'h00C7D713;
    mem['h0223] <= 32'h01479793;
    mem['h0224] <= 32'h00E7E7B3;
    mem['h0225] <= 32'hF2F42423;
    mem['h0226] <= 32'hF1842703;
    mem['h0227] <= 32'hF2842783;
    mem['h0228] <= 32'h00F70733;
    mem['h0229] <= 32'hFEC42783;
    mem['h022A] <= 32'h00479793;
    mem['h022B] <= 32'hFF078793;
    mem['h022C] <= 32'h008787B3;
    mem['h022D] <= 32'hF637C783;
    mem['h022E] <= 32'h00279793;
    mem['h022F] <= 32'hFF078793;
    mem['h0230] <= 32'h008787B3;
    mem['h0231] <= 32'hEDC7A783;
    mem['h0232] <= 32'h00F707B3;
    mem['h0233] <= 32'hF0F42C23;
    mem['h0234] <= 32'hF4842703;
    mem['h0235] <= 32'hF1842783;
    mem['h0236] <= 32'h00F747B3;
    mem['h0237] <= 32'h0087D713;
    mem['h0238] <= 32'h01879793;
    mem['h0239] <= 32'h00E7E7B3;
    mem['h023A] <= 32'hF4F42423;
    mem['h023B] <= 32'hF3842703;
    mem['h023C] <= 32'hF4842783;
    mem['h023D] <= 32'h00F707B3;
    mem['h023E] <= 32'hF2F42C23;
    mem['h023F] <= 32'hF2842703;
    mem['h0240] <= 32'hF3842783;
    mem['h0241] <= 32'h00F747B3;
    mem['h0242] <= 32'h0077D713;
    mem['h0243] <= 32'h01979793;
    mem['h0244] <= 32'h00E7E7B3;
    mem['h0245] <= 32'hF2F42423;
    mem['h0246] <= 32'hF0C42703;
    mem['h0247] <= 32'hF2042783;
    mem['h0248] <= 32'h00F70733;
    mem['h0249] <= 32'hFEC42783;
    mem['h024A] <= 32'h00479793;
    mem['h024B] <= 32'hFF078793;
    mem['h024C] <= 32'h008787B3;
    mem['h024D] <= 32'hF647C783;
    mem['h024E] <= 32'h00279793;
    mem['h024F] <= 32'hFF078793;
    mem['h0250] <= 32'h008787B3;
    mem['h0251] <= 32'hEDC7A783;
    mem['h0252] <= 32'h00F707B3;
    mem['h0253] <= 32'hF0F42623;
    mem['h0254] <= 32'hF4842703;
    mem['h0255] <= 32'hF0C42783;
    mem['h0256] <= 32'h00F747B3;
    mem['h0257] <= 32'h01079713;
    mem['h0258] <= 32'h0107D793;
    mem['h0259] <= 32'h00E7E7B3;
    mem['h025A] <= 32'hF4F42423;
    mem['h025B] <= 32'hF3442703;
    mem['h025C] <= 32'hF4842783;
    mem['h025D] <= 32'h00F707B3;
    mem['h025E] <= 32'hF2F42A23;
    mem['h025F] <= 32'hF2042703;
    mem['h0260] <= 32'hF3442783;
    mem['h0261] <= 32'h00F747B3;
    mem['h0262] <= 32'h00C7D713;
    mem['h0263] <= 32'h01479793;
    mem['h0264] <= 32'h00E7E7B3;
    mem['h0265] <= 32'hF2F42023;
    mem['h0266] <= 32'hF0C42703;
    mem['h0267] <= 32'hF2042783;
    mem['h0268] <= 32'h00F70733;
    mem['h0269] <= 32'hFEC42783;
    mem['h026A] <= 32'h00479793;
    mem['h026B] <= 32'hFF078793;
    mem['h026C] <= 32'h008787B3;
    mem['h026D] <= 32'hF657C783;
    mem['h026E] <= 32'h00279793;
    mem['h026F] <= 32'hFF078793;
    mem['h0270] <= 32'h008787B3;
    mem['h0271] <= 32'hEDC7A783;
    mem['h0272] <= 32'h00F707B3;
    mem['h0273] <= 32'hF0F42623;
    mem['h0274] <= 32'hF4842703;
    mem['h0275] <= 32'hF0C42783;
    mem['h0276] <= 32'h00F747B3;
    mem['h0277] <= 32'h0087D713;
    mem['h0278] <= 32'h01879793;
    mem['h0279] <= 32'h00E7E7B3;
    mem['h027A] <= 32'hF4F42423;
    mem['h027B] <= 32'hF3442703;
    mem['h027C] <= 32'hF4842783;
    mem['h027D] <= 32'h00F707B3;
    mem['h027E] <= 32'hF2F42A23;
    mem['h027F] <= 32'hF2042703;
    mem['h0280] <= 32'hF3442783;
    mem['h0281] <= 32'h00F747B3;
    mem['h0282] <= 32'h0077D713;
    mem['h0283] <= 32'h01979793;
    mem['h0284] <= 32'h00E7E7B3;
    mem['h0285] <= 32'hF2F42023;
    mem['h0286] <= 32'hF1042703;
    mem['h0287] <= 32'hF2442783;
    mem['h0288] <= 32'h00F70733;
    mem['h0289] <= 32'hFEC42783;
    mem['h028A] <= 32'h00479793;
    mem['h028B] <= 32'hFF078793;
    mem['h028C] <= 32'h008787B3;
    mem['h028D] <= 32'hF667C783;
    mem['h028E] <= 32'h00279793;
    mem['h028F] <= 32'hFF078793;
    mem['h0290] <= 32'h008787B3;
    mem['h0291] <= 32'hEDC7A783;
    mem['h0292] <= 32'h00F707B3;
    mem['h0293] <= 32'hF0F42823;
    mem['h0294] <= 32'hF3C42703;
    mem['h0295] <= 32'hF1042783;
    mem['h0296] <= 32'h00F747B3;
    mem['h0297] <= 32'h01079713;
    mem['h0298] <= 32'h0107D793;
    mem['h0299] <= 32'h00E7E7B3;
    mem['h029A] <= 32'hF2F42E23;
    mem['h029B] <= 32'hF3842703;
    mem['h029C] <= 32'hF3C42783;
    mem['h029D] <= 32'h00F707B3;
    mem['h029E] <= 32'hF2F42C23;
    mem['h029F] <= 32'hF2442703;
    mem['h02A0] <= 32'hF3842783;
    mem['h02A1] <= 32'h00F747B3;
    mem['h02A2] <= 32'h00C7D713;
    mem['h02A3] <= 32'h01479793;
    mem['h02A4] <= 32'h00E7E7B3;
    mem['h02A5] <= 32'hF2F42223;
    mem['h02A6] <= 32'hF1042703;
    mem['h02A7] <= 32'hF2442783;
    mem['h02A8] <= 32'h00F70733;
    mem['h02A9] <= 32'hFEC42783;
    mem['h02AA] <= 32'h00479793;
    mem['h02AB] <= 32'hFF078793;
    mem['h02AC] <= 32'h008787B3;
    mem['h02AD] <= 32'hF677C783;
    mem['h02AE] <= 32'h00279793;
    mem['h02AF] <= 32'hFF078793;
    mem['h02B0] <= 32'h008787B3;
    mem['h02B1] <= 32'hEDC7A783;
    mem['h02B2] <= 32'h00F707B3;
    mem['h02B3] <= 32'hF0F42823;
    mem['h02B4] <= 32'hF3C42703;
    mem['h02B5] <= 32'hF1042783;
    mem['h02B6] <= 32'h00F747B3;
    mem['h02B7] <= 32'h0087D713;
    mem['h02B8] <= 32'h01879793;
    mem['h02B9] <= 32'h00E7E7B3;
    mem['h02BA] <= 32'hF2F42E23;
    mem['h02BB] <= 32'hF3842703;
    mem['h02BC] <= 32'hF3C42783;
    mem['h02BD] <= 32'h00F707B3;
    mem['h02BE] <= 32'hF2F42C23;
    mem['h02BF] <= 32'hF2442703;
    mem['h02C0] <= 32'hF3842783;
    mem['h02C1] <= 32'h00F747B3;
    mem['h02C2] <= 32'h0077D713;
    mem['h02C3] <= 32'h01979793;
    mem['h02C4] <= 32'h00E7E7B3;
    mem['h02C5] <= 32'hF2F42223;
    mem['h02C6] <= 32'hF1442703;
    mem['h02C7] <= 32'hF2842783;
    mem['h02C8] <= 32'h00F70733;
    mem['h02C9] <= 32'hFEC42783;
    mem['h02CA] <= 32'h00479793;
    mem['h02CB] <= 32'hFF078793;
    mem['h02CC] <= 32'h008787B3;
    mem['h02CD] <= 32'hF687C783;
    mem['h02CE] <= 32'h00279793;
    mem['h02CF] <= 32'hFF078793;
    mem['h02D0] <= 32'h008787B3;
    mem['h02D1] <= 32'hEDC7A783;
    mem['h02D2] <= 32'h00F707B3;
    mem['h02D3] <= 32'hF0F42A23;
    mem['h02D4] <= 32'hF4042703;
    mem['h02D5] <= 32'hF1442783;
    mem['h02D6] <= 32'h00F747B3;
    mem['h02D7] <= 32'h01079713;
    mem['h02D8] <= 32'h0107D793;
    mem['h02D9] <= 32'h00E7E7B3;
    mem['h02DA] <= 32'hF4F42023;
    mem['h02DB] <= 32'hF2C42703;
    mem['h02DC] <= 32'hF4042783;
    mem['h02DD] <= 32'h00F707B3;
    mem['h02DE] <= 32'hF2F42623;
    mem['h02DF] <= 32'hF2842703;
    mem['h02E0] <= 32'hF2C42783;
    mem['h02E1] <= 32'h00F747B3;
    mem['h02E2] <= 32'h00C7D713;
    mem['h02E3] <= 32'h01479793;
    mem['h02E4] <= 32'h00E7E7B3;
    mem['h02E5] <= 32'hF2F42423;
    mem['h02E6] <= 32'hF1442703;
    mem['h02E7] <= 32'hF2842783;
    mem['h02E8] <= 32'h00F70733;
    mem['h02E9] <= 32'hFEC42783;
    mem['h02EA] <= 32'h00479793;
    mem['h02EB] <= 32'hFF078793;
    mem['h02EC] <= 32'h008787B3;
    mem['h02ED] <= 32'hF697C783;
    mem['h02EE] <= 32'h00279793;
    mem['h02EF] <= 32'hFF078793;
    mem['h02F0] <= 32'h008787B3;
    mem['h02F1] <= 32'hEDC7A783;
    mem['h02F2] <= 32'h00F707B3;
    mem['h02F3] <= 32'hF0F42A23;
    mem['h02F4] <= 32'hF4042703;
    mem['h02F5] <= 32'hF1442783;
    mem['h02F6] <= 32'h00F747B3;
    mem['h02F7] <= 32'h0087D713;
    mem['h02F8] <= 32'h01879793;
    mem['h02F9] <= 32'h00E7E7B3;
    mem['h02FA] <= 32'hF4F42023;
    mem['h02FB] <= 32'hF2C42703;
    mem['h02FC] <= 32'hF4042783;
    mem['h02FD] <= 32'h00F707B3;
    mem['h02FE] <= 32'hF2F42623;
    mem['h02FF] <= 32'hF2842703;
    mem['h0300] <= 32'hF2C42783;
    mem['h0301] <= 32'h00F747B3;
    mem['h0302] <= 32'h0077D713;
    mem['h0303] <= 32'h01979793;
    mem['h0304] <= 32'h00E7E7B3;
    mem['h0305] <= 32'hF2F42423;
    mem['h0306] <= 32'hF1842703;
    mem['h0307] <= 32'hF1C42783;
    mem['h0308] <= 32'h00F70733;
    mem['h0309] <= 32'hFEC42783;
    mem['h030A] <= 32'h00479793;
    mem['h030B] <= 32'hFF078793;
    mem['h030C] <= 32'h008787B3;
    mem['h030D] <= 32'hF6A7C783;
    mem['h030E] <= 32'h00279793;
    mem['h030F] <= 32'hFF078793;
    mem['h0310] <= 32'h008787B3;
    mem['h0311] <= 32'hEDC7A783;
    mem['h0312] <= 32'h00F707B3;
    mem['h0313] <= 32'hF0F42C23;
    mem['h0314] <= 32'hF4442703;
    mem['h0315] <= 32'hF1842783;
    mem['h0316] <= 32'h00F747B3;
    mem['h0317] <= 32'h01079713;
    mem['h0318] <= 32'h0107D793;
    mem['h0319] <= 32'h00E7E7B3;
    mem['h031A] <= 32'hF4F42223;
    mem['h031B] <= 32'hF3042703;
    mem['h031C] <= 32'hF4442783;
    mem['h031D] <= 32'h00F707B3;
    mem['h031E] <= 32'hF2F42823;
    mem['h031F] <= 32'hF1C42703;
    mem['h0320] <= 32'hF3042783;
    mem['h0321] <= 32'h00F747B3;
    mem['h0322] <= 32'h00C7D713;
    mem['h0323] <= 32'h01479793;
    mem['h0324] <= 32'h00E7E7B3;
    mem['h0325] <= 32'hF0F42E23;
    mem['h0326] <= 32'hF1842703;
    mem['h0327] <= 32'hF1C42783;
    mem['h0328] <= 32'h00F70733;
    mem['h0329] <= 32'hFEC42783;
    mem['h032A] <= 32'h00479793;
    mem['h032B] <= 32'hFF078793;
    mem['h032C] <= 32'h008787B3;
    mem['h032D] <= 32'hF6B7C783;
    mem['h032E] <= 32'h00279793;
    mem['h032F] <= 32'hFF078793;
    mem['h0330] <= 32'h008787B3;
    mem['h0331] <= 32'hEDC7A783;
    mem['h0332] <= 32'h00F707B3;
    mem['h0333] <= 32'hF0F42C23;
    mem['h0334] <= 32'hF4442703;
    mem['h0335] <= 32'hF1842783;
    mem['h0336] <= 32'h00F747B3;
    mem['h0337] <= 32'h0087D713;
    mem['h0338] <= 32'h01879793;
    mem['h0339] <= 32'h00E7E7B3;
    mem['h033A] <= 32'hF4F42223;
    mem['h033B] <= 32'hF3042703;
    mem['h033C] <= 32'hF4442783;
    mem['h033D] <= 32'h00F707B3;
    mem['h033E] <= 32'hF2F42823;
    mem['h033F] <= 32'hF1C42703;
    mem['h0340] <= 32'hF3042783;
    mem['h0341] <= 32'h00F747B3;
    mem['h0342] <= 32'h0077D713;
    mem['h0343] <= 32'h01979793;
    mem['h0344] <= 32'h00E7E7B3;
    mem['h0345] <= 32'hF0F42E23;
    mem['h0346] <= 32'hFEC42783;
    mem['h0347] <= 32'h00178793;
    mem['h0348] <= 32'hFEF42623;
    mem['h0349] <= 32'hFEC42703;
    mem['h034A] <= 32'h00900793;
    mem['h034B] <= 32'hFEE7D663;
    mem['h034C] <= 32'hFE042623;
    mem['h034D] <= 32'h0740006F;
    mem['h034E] <= 32'hEBC42703;
    mem['h034F] <= 32'hFEC42783;
    mem['h0350] <= 32'h01078793;
    mem['h0351] <= 32'h00279793;
    mem['h0352] <= 32'h00F707B3;
    mem['h0353] <= 32'h0007A703;
    mem['h0354] <= 32'hFEC42783;
    mem['h0355] <= 32'h00279793;
    mem['h0356] <= 32'hFF078793;
    mem['h0357] <= 32'h008787B3;
    mem['h0358] <= 32'hF1C7A683;
    mem['h0359] <= 32'hFEC42783;
    mem['h035A] <= 32'h00878793;
    mem['h035B] <= 32'h00279793;
    mem['h035C] <= 32'hFF078793;
    mem['h035D] <= 32'h008787B3;
    mem['h035E] <= 32'hF1C7A783;
    mem['h035F] <= 32'h00F6C7B3;
    mem['h0360] <= 32'h00F74733;
    mem['h0361] <= 32'hEBC42683;
    mem['h0362] <= 32'hFEC42783;
    mem['h0363] <= 32'h01078793;
    mem['h0364] <= 32'h00279793;
    mem['h0365] <= 32'h00F687B3;
    mem['h0366] <= 32'h00E7A023;
    mem['h0367] <= 32'hFEC42783;
    mem['h0368] <= 32'h00178793;
    mem['h0369] <= 32'hFEF42623;
    mem['h036A] <= 32'hFEC42703;
    mem['h036B] <= 32'h00700793;
    mem['h036C] <= 32'hF8E7D4E3;
    mem['h036D] <= 32'h00000013;
    mem['h036E] <= 32'h00000013;
    mem['h036F] <= 32'h14C12083;
    mem['h0370] <= 32'h14812403;
    mem['h0371] <= 32'h15010113;
    mem['h0372] <= 32'h00008067;
    mem['h0373] <= 32'hFD010113;
    mem['h0374] <= 32'h02112623;
    mem['h0375] <= 32'h02812423;
    mem['h0376] <= 32'h03010413;
    mem['h0377] <= 32'hFCA42E23;
    mem['h0378] <= 32'hFCB42C23;
    mem['h0379] <= 32'hFCC42A23;
    mem['h037A] <= 32'hFCD42823;
    mem['h037B] <= 32'hFD842783;
    mem['h037C] <= 32'h00078E63;
    mem['h037D] <= 32'hFD842703;
    mem['h037E] <= 32'h02000793;
    mem['h037F] <= 32'h00E7E863;
    mem['h0380] <= 32'hFD042703;
    mem['h0381] <= 32'h02000793;
    mem['h0382] <= 32'h00E7F663;
    mem['h0383] <= 32'hFFF00793;
    mem['h0384] <= 32'h1000006F;
    mem['h0385] <= 32'hFE042623;
    mem['h0386] <= 32'h0400006F;
    mem['h0387] <= 32'h001017B7;
    mem['h0388] <= 32'h39878713;
    mem['h0389] <= 32'hFEC42783;
    mem['h038A] <= 32'h00279793;
    mem['h038B] <= 32'h00F707B3;
    mem['h038C] <= 32'h0007A703;
    mem['h038D] <= 32'hFDC42683;
    mem['h038E] <= 32'hFEC42783;
    mem['h038F] <= 32'h01078793;
    mem['h0390] <= 32'h00279793;
    mem['h0391] <= 32'h00F687B3;
    mem['h0392] <= 32'h00E7A023;
    mem['h0393] <= 32'hFEC42783;
    mem['h0394] <= 32'h00178793;
    mem['h0395] <= 32'hFEF42623;
    mem['h0396] <= 32'hFEC42703;
    mem['h0397] <= 32'h00700793;
    mem['h0398] <= 32'hFAE7FEE3;
    mem['h0399] <= 32'hFDC42783;
    mem['h039A] <= 32'h0407A703;
    mem['h039B] <= 32'hFD042783;
    mem['h039C] <= 32'h00879693;
    mem['h039D] <= 32'hFD842783;
    mem['h039E] <= 32'h00F6C7B3;
    mem['h039F] <= 32'h00F74733;
    mem['h03A0] <= 32'h010107B7;
    mem['h03A1] <= 32'h00F74733;
    mem['h03A2] <= 32'hFDC42783;
    mem['h03A3] <= 32'h04E7A023;
    mem['h03A4] <= 32'hFDC42783;
    mem['h03A5] <= 32'h0607A023;
    mem['h03A6] <= 32'hFDC42783;
    mem['h03A7] <= 32'h0607A223;
    mem['h03A8] <= 32'hFDC42783;
    mem['h03A9] <= 32'h0607A423;
    mem['h03AA] <= 32'hFDC42783;
    mem['h03AB] <= 32'hFD842703;
    mem['h03AC] <= 32'h06E7A623;
    mem['h03AD] <= 32'hFD042783;
    mem['h03AE] <= 32'hFEF42623;
    mem['h03AF] <= 32'h0200006F;
    mem['h03B0] <= 32'hFDC42703;
    mem['h03B1] <= 32'hFEC42783;
    mem['h03B2] <= 32'h00F707B3;
    mem['h03B3] <= 32'h00078023;
    mem['h03B4] <= 32'hFEC42783;
    mem['h03B5] <= 32'h00178793;
    mem['h03B6] <= 32'hFEF42623;
    mem['h03B7] <= 32'hFEC42703;
    mem['h03B8] <= 32'h03F00793;
    mem['h03B9] <= 32'hFCE7FEE3;
    mem['h03BA] <= 32'hFD042783;
    mem['h03BB] <= 32'h02078063;
    mem['h03BC] <= 32'hFD042603;
    mem['h03BD] <= 32'hFD442583;
    mem['h03BE] <= 32'hFDC42503;
    mem['h03BF] <= 32'h028000EF;
    mem['h03C0] <= 32'hFDC42783;
    mem['h03C1] <= 32'h04000713;
    mem['h03C2] <= 32'h06E7A423;
    mem['h03C3] <= 32'h00000793;
    mem['h03C4] <= 32'h00078513;
    mem['h03C5] <= 32'h02C12083;
    mem['h03C6] <= 32'h02812403;
    mem['h03C7] <= 32'h03010113;
    mem['h03C8] <= 32'h00008067;
    mem['h03C9] <= 32'hFD010113;
    mem['h03CA] <= 32'h02112623;
    mem['h03CB] <= 32'h02812423;
    mem['h03CC] <= 32'h03010413;
    mem['h03CD] <= 32'hFCA42E23;
    mem['h03CE] <= 32'hFCB42C23;
    mem['h03CF] <= 32'hFCC42A23;
    mem['h03D0] <= 32'hFE042623;
    mem['h03D1] <= 32'h0A80006F;
    mem['h03D2] <= 32'hFDC42783;
    mem['h03D3] <= 32'h0687A703;
    mem['h03D4] <= 32'h04000793;
    mem['h03D5] <= 32'h04F71E63;
    mem['h03D6] <= 32'hFDC42783;
    mem['h03D7] <= 32'h0607A703;
    mem['h03D8] <= 32'hFDC42783;
    mem['h03D9] <= 32'h0687A783;
    mem['h03DA] <= 32'h00F70733;
    mem['h03DB] <= 32'hFDC42783;
    mem['h03DC] <= 32'h06E7A023;
    mem['h03DD] <= 32'hFDC42783;
    mem['h03DE] <= 32'h0607A703;
    mem['h03DF] <= 32'hFDC42783;
    mem['h03E0] <= 32'h0687A783;
    mem['h03E1] <= 32'h00F77C63;
    mem['h03E2] <= 32'hFDC42783;
    mem['h03E3] <= 32'h0647A783;
    mem['h03E4] <= 32'h00178713;
    mem['h03E5] <= 32'hFDC42783;
    mem['h03E6] <= 32'h06E7A223;
    mem['h03E7] <= 32'h00000593;
    mem['h03E8] <= 32'hFDC42503;
    mem['h03E9] <= 32'hBCCFF0EF;
    mem['h03EA] <= 32'hFDC42783;
    mem['h03EB] <= 32'h0607A423;
    mem['h03EC] <= 32'hFD842703;
    mem['h03ED] <= 32'hFEC42783;
    mem['h03EE] <= 32'h00F70733;
    mem['h03EF] <= 32'hFDC42783;
    mem['h03F0] <= 32'h0687A783;
    mem['h03F1] <= 32'h00178613;
    mem['h03F2] <= 32'hFDC42683;
    mem['h03F3] <= 32'h06C6A423;
    mem['h03F4] <= 32'h00074703;
    mem['h03F5] <= 32'hFDC42683;
    mem['h03F6] <= 32'h00F687B3;
    mem['h03F7] <= 32'h00E78023;
    mem['h03F8] <= 32'hFEC42783;
    mem['h03F9] <= 32'h00178793;
    mem['h03FA] <= 32'hFEF42623;
    mem['h03FB] <= 32'hFEC42703;
    mem['h03FC] <= 32'hFD442783;
    mem['h03FD] <= 32'hF4F76AE3;
    mem['h03FE] <= 32'h00000013;
    mem['h03FF] <= 32'h00000013;
    mem['h0400] <= 32'h02C12083;
    mem['h0401] <= 32'h02812403;
    mem['h0402] <= 32'h03010113;
    mem['h0403] <= 32'h00008067;
    mem['h0404] <= 32'hFD010113;
    mem['h0405] <= 32'h02112623;
    mem['h0406] <= 32'h02812423;
    mem['h0407] <= 32'h03010413;
    mem['h0408] <= 32'hFCA42E23;
    mem['h0409] <= 32'hFCB42C23;
    mem['h040A] <= 32'hFDC42783;
    mem['h040B] <= 32'h0607A703;
    mem['h040C] <= 32'hFDC42783;
    mem['h040D] <= 32'h0687A783;
    mem['h040E] <= 32'h00F70733;
    mem['h040F] <= 32'hFDC42783;
    mem['h0410] <= 32'h06E7A023;
    mem['h0411] <= 32'hFDC42783;
    mem['h0412] <= 32'h0607A703;
    mem['h0413] <= 32'hFDC42783;
    mem['h0414] <= 32'h0687A783;
    mem['h0415] <= 32'h02F77E63;
    mem['h0416] <= 32'hFDC42783;
    mem['h0417] <= 32'h0647A783;
    mem['h0418] <= 32'h00178713;
    mem['h0419] <= 32'hFDC42783;
    mem['h041A] <= 32'h06E7A223;
    mem['h041B] <= 32'h0240006F;
    mem['h041C] <= 32'hFDC42783;
    mem['h041D] <= 32'h0687A783;
    mem['h041E] <= 32'h00178693;
    mem['h041F] <= 32'hFDC42703;
    mem['h0420] <= 32'h06D72423;
    mem['h0421] <= 32'hFDC42703;
    mem['h0422] <= 32'h00F707B3;
    mem['h0423] <= 32'h00078023;
    mem['h0424] <= 32'hFDC42783;
    mem['h0425] <= 32'h0687A703;
    mem['h0426] <= 32'h03F00793;
    mem['h0427] <= 32'hFCE7FAE3;
    mem['h0428] <= 32'h00100593;
    mem['h0429] <= 32'hFDC42503;
    mem['h042A] <= 32'hAC8FF0EF;
    mem['h042B] <= 32'hFE042623;
    mem['h042C] <= 32'h0500006F;
    mem['h042D] <= 32'hFEC42783;
    mem['h042E] <= 32'h0027D793;
    mem['h042F] <= 32'hFDC42703;
    mem['h0430] <= 32'h01078793;
    mem['h0431] <= 32'h00279793;
    mem['h0432] <= 32'h00F707B3;
    mem['h0433] <= 32'h0007A703;
    mem['h0434] <= 32'hFEC42783;
    mem['h0435] <= 32'h0037F793;
    mem['h0436] <= 32'h00379793;
    mem['h0437] <= 32'h00F756B3;
    mem['h0438] <= 32'hFD842703;
    mem['h0439] <= 32'hFEC42783;
    mem['h043A] <= 32'h00F707B3;
    mem['h043B] <= 32'h0FF6F713;
    mem['h043C] <= 32'h00E78023;
    mem['h043D] <= 32'hFEC42783;
    mem['h043E] <= 32'h00178793;
    mem['h043F] <= 32'hFEF42623;
    mem['h0440] <= 32'hFDC42783;
    mem['h0441] <= 32'h06C7A783;
    mem['h0442] <= 32'hFEC42703;
    mem['h0443] <= 32'hFAF764E3;
    mem['h0444] <= 32'h00000013;
    mem['h0445] <= 32'h00000013;
    mem['h0446] <= 32'h02C12083;
    mem['h0447] <= 32'h02812403;
    mem['h0448] <= 32'h03010113;
    mem['h0449] <= 32'h00008067;
    mem['h044A] <= 32'hF6010113;
    mem['h044B] <= 32'h08112E23;
    mem['h044C] <= 32'h08812C23;
    mem['h044D] <= 32'h0A010413;
    mem['h044E] <= 32'hF6A42E23;
    mem['h044F] <= 32'hF6B42C23;
    mem['h0450] <= 32'hF6C42A23;
    mem['h0451] <= 32'hF6D42823;
    mem['h0452] <= 32'hF6E42623;
    mem['h0453] <= 32'hF6F42423;
    mem['h0454] <= 32'hF8040793;
    mem['h0455] <= 32'hF7042683;
    mem['h0456] <= 32'hF7442603;
    mem['h0457] <= 32'hF7842583;
    mem['h0458] <= 32'h00078513;
    mem['h0459] <= 32'hC69FF0EF;
    mem['h045A] <= 32'h00050793;
    mem['h045B] <= 32'h00078663;
    mem['h045C] <= 32'hFFF00793;
    mem['h045D] <= 32'h02C0006F;
    mem['h045E] <= 32'hF8040793;
    mem['h045F] <= 32'hF6842603;
    mem['h0460] <= 32'hF6C42583;
    mem['h0461] <= 32'h00078513;
    mem['h0462] <= 32'hD9DFF0EF;
    mem['h0463] <= 32'hF8040793;
    mem['h0464] <= 32'hF7C42583;
    mem['h0465] <= 32'h00078513;
    mem['h0466] <= 32'hE79FF0EF;
    mem['h0467] <= 32'h00000793;
    mem['h0468] <= 32'h00078513;
    mem['h0469] <= 32'h09C12083;
    mem['h046A] <= 32'h09812403;
    mem['h046B] <= 32'h0A010113;
    mem['h046C] <= 32'h00008067;
    mem['h046D] <= 32'hFD010113;
    mem['h046E] <= 32'h02812623;
    mem['h046F] <= 32'h03010413;
    mem['h0470] <= 32'hFCA42E23;
    mem['h0471] <= 32'hFCB42C23;
    mem['h0472] <= 32'hFCC42A23;
    mem['h0473] <= 32'hFDC42783;
    mem['h0474] <= 32'hFEF42423;
    mem['h0475] <= 32'hFD842783;
    mem['h0476] <= 32'hFEF403A3;
    mem['h0477] <= 32'hFE042623;
    mem['h0478] <= 32'h0240006F;
    mem['h0479] <= 32'hFE842703;
    mem['h047A] <= 32'hFEC42783;
    mem['h047B] <= 32'h00F707B3;
    mem['h047C] <= 32'hFE744703;
    mem['h047D] <= 32'h00E78023;
    mem['h047E] <= 32'hFEC42783;
    mem['h047F] <= 32'h00178793;
    mem['h0480] <= 32'hFEF42623;
    mem['h0481] <= 32'hFEC42703;
    mem['h0482] <= 32'hFD442783;
    mem['h0483] <= 32'hFCF76CE3;
    mem['h0484] <= 32'hFDC42783;
    mem['h0485] <= 32'h00078513;
    mem['h0486] <= 32'h02C12403;
    mem['h0487] <= 32'h03010113;
    mem['h0488] <= 32'h00008067;
    mem['h0489] <= 32'hFD010113;
    mem['h048A] <= 32'h02812623;
    mem['h048B] <= 32'h03010413;
    mem['h048C] <= 32'hFCA42E23;
    mem['h048D] <= 32'hFCB42C23;
    mem['h048E] <= 32'hFCC42A23;
    mem['h048F] <= 32'hFDC42783;
    mem['h0490] <= 32'hFEF42423;
    mem['h0491] <= 32'hFD842783;
    mem['h0492] <= 32'hFEF42223;
    mem['h0493] <= 32'hFE042623;
    mem['h0494] <= 32'h0300006F;
    mem['h0495] <= 32'hFE442703;
    mem['h0496] <= 32'hFEC42783;
    mem['h0497] <= 32'h00F70733;
    mem['h0498] <= 32'hFE842683;
    mem['h0499] <= 32'hFEC42783;
    mem['h049A] <= 32'h00F687B3;
    mem['h049B] <= 32'h00074703;
    mem['h049C] <= 32'h00E78023;
    mem['h049D] <= 32'hFEC42783;
    mem['h049E] <= 32'h00178793;
    mem['h049F] <= 32'hFEF42623;
    mem['h04A0] <= 32'hFEC42703;
    mem['h04A1] <= 32'hFD442783;
    mem['h04A2] <= 32'hFCF766E3;
    mem['h04A3] <= 32'hFDC42783;
    mem['h04A4] <= 32'h00078513;
    mem['h04A5] <= 32'h02C12403;
    mem['h04A6] <= 32'h03010113;
    mem['h04A7] <= 32'h00008067;
    mem['h04A8] <= 32'hFD010113;
    mem['h04A9] <= 32'h02812623;
    mem['h04AA] <= 32'h03010413;
    mem['h04AB] <= 32'hFCA42E23;
    mem['h04AC] <= 32'hFCB42C23;
    mem['h04AD] <= 32'hFCC42A23;
    mem['h04AE] <= 32'hFDC42783;
    mem['h04AF] <= 32'hFEF42423;
    mem['h04B0] <= 32'hFD842783;
    mem['h04B1] <= 32'hFEF42223;
    mem['h04B2] <= 32'hFE042623;
    mem['h04B3] <= 32'h0600006F;
    mem['h04B4] <= 32'hFE842703;
    mem['h04B5] <= 32'hFEC42783;
    mem['h04B6] <= 32'h00F707B3;
    mem['h04B7] <= 32'h0007C703;
    mem['h04B8] <= 32'hFE442683;
    mem['h04B9] <= 32'hFEC42783;
    mem['h04BA] <= 32'h00F687B3;
    mem['h04BB] <= 32'h0007C783;
    mem['h04BC] <= 32'h02F70863;
    mem['h04BD] <= 32'hFE842703;
    mem['h04BE] <= 32'hFEC42783;
    mem['h04BF] <= 32'h00F707B3;
    mem['h04C0] <= 32'h0007C783;
    mem['h04C1] <= 32'h00078693;
    mem['h04C2] <= 32'hFE442703;
    mem['h04C3] <= 32'hFEC42783;
    mem['h04C4] <= 32'h00F707B3;
    mem['h04C5] <= 32'h0007C783;
    mem['h04C6] <= 32'h40F687B3;
    mem['h04C7] <= 32'h0200006F;
    mem['h04C8] <= 32'hFEC42783;
    mem['h04C9] <= 32'h00178793;
    mem['h04CA] <= 32'hFEF42623;
    mem['h04CB] <= 32'hFEC42703;
    mem['h04CC] <= 32'hFD442783;
    mem['h04CD] <= 32'hF8F76EE3;
    mem['h04CE] <= 32'h00000793;
    mem['h04CF] <= 32'h00078513;
    mem['h04D0] <= 32'h02C12403;
    mem['h04D1] <= 32'h03010113;
    mem['h04D2] <= 32'h00008067;
    mem['h04D3] <= 32'hFD010113;
    mem['h04D4] <= 32'h02812623;
    mem['h04D5] <= 32'h03010413;
    mem['h04D6] <= 32'hFCA42E23;
    mem['h04D7] <= 32'hFE042623;
    mem['h04D8] <= 32'h0100006F;
    mem['h04D9] <= 32'hFEC42783;
    mem['h04DA] <= 32'h00178793;
    mem['h04DB] <= 32'hFEF42623;
    mem['h04DC] <= 32'hFDC42703;
    mem['h04DD] <= 32'hFEC42783;
    mem['h04DE] <= 32'h00F707B3;
    mem['h04DF] <= 32'h0007C783;
    mem['h04E0] <= 32'hFE0792E3;
    mem['h04E1] <= 32'hFEC42783;
    mem['h04E2] <= 32'h00078513;
    mem['h04E3] <= 32'h02C12403;
    mem['h04E4] <= 32'h03010113;
    mem['h04E5] <= 32'h00008067;
    mem['h04E6] <= 32'h6A09E667;
    mem['h04E7] <= 32'hBB67AE85;
    mem['h04E8] <= 32'h3C6EF372;
    mem['h04E9] <= 32'hA54FF53A;
    mem['h04EA] <= 32'h510E527F;
    mem['h04EB] <= 32'h9B05688C;
    mem['h04EC] <= 32'h1F83D9AB;
    mem['h04ED] <= 32'h5BE0CD19;
    mem['h04EE] <= 32'h03020100;
    mem['h04EF] <= 32'h07060504;
    mem['h04F0] <= 32'h0B0A0908;
    mem['h04F1] <= 32'h0F0E0D0C;
    mem['h04F2] <= 32'h08040A0E;
    mem['h04F3] <= 32'h060D0F09;
    mem['h04F4] <= 32'h02000C01;
    mem['h04F5] <= 32'h0305070B;
    mem['h04F6] <= 32'h000C080B;
    mem['h04F7] <= 32'h0D0F0205;
    mem['h04F8] <= 32'h06030E0A;
    mem['h04F9] <= 32'h04090107;
    mem['h04FA] <= 32'h01030907;
    mem['h04FB] <= 32'h0E0B0C0D;
    mem['h04FC] <= 32'h0A050602;
    mem['h04FD] <= 32'h080F0004;
    mem['h04FE] <= 32'h07050009;
    mem['h04FF] <= 32'h0F0A0402;
    mem['h0500] <= 32'h0C0B010E;
    mem['h0501] <= 32'h0D030806;
    mem['h0502] <= 32'h0A060C02;
    mem['h0503] <= 32'h03080B00;
    mem['h0504] <= 32'h05070D04;
    mem['h0505] <= 32'h09010E0F;
    mem['h0506] <= 32'h0F01050C;
    mem['h0507] <= 32'h0A040D0E;
    mem['h0508] <= 32'h03060700;
    mem['h0509] <= 32'h0B080209;
    mem['h050A] <= 32'h0E070B0D;
    mem['h050B] <= 32'h0903010C;
    mem['h050C] <= 32'h040F0005;
    mem['h050D] <= 32'h0A020608;
    mem['h050E] <= 32'h090E0F06;
    mem['h050F] <= 32'h0800030B;
    mem['h0510] <= 32'h070D020C;
    mem['h0511] <= 32'h050A0401;
    mem['h0512] <= 32'h0408020A;
    mem['h0513] <= 32'h05010607;
    mem['h0514] <= 32'h0E090B0F;
    mem['h0515] <= 32'h000D0C03;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

  always @(posedge clk) begin
    if (wen) mem[waddr] <= wdata;
  end

endmodule
