-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.20810055865921787, 0.5921787709497207, 0.9762569832402235]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_3CLK_087b5579 is
port(
 clk : in std_logic;
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_3CLK_087b5579;
architecture arch of uint320_mul_3CLK_087b5579 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 3;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
-- Stage 1
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
-- Stage 2
signal REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
signal COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_2a7e]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8597]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_fec3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_09f7]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4c9a]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_b459]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_d7df]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_475c]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_958d]
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_fe6a]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_0a85]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_9973]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_0285]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_de17]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_ee02]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_1838]
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_83f1]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_42fd]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_866a]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_9e29]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_3e3b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_0a27]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_33f6]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_886b]
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204]
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3]
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_c44d]
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_9ca18c4f port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_41a2906e port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_eec62983 port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right,
FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285 : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_1CLK_9324e8e6 port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0f464748 port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right,
FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_1CLK_ec635a74 port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1 : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_0320092f port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right,
FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right,
FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204 : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : 0 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output);

-- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d : 1 clocks latency
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d : entity work.BIN_OP_PLUS_uint64_t_uint64_t_1CLK_8f2211ba port map (
clk,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right,
FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- Registers
 -- Stage 0
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 -- Stage 1
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left,
 -- Stage 2
 REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output,
 FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_7dfc_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_7dfc_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_7dfc_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_7dfc_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_e477_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_7dfc_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_7a4b_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_123a_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_e477_DUPLICATE_632a_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_e477_DUPLICATE_226e_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_acaf_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_5233_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse := to_unsigned(0, 64);
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_7dfc] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_7dfc_return_output := u320_t_NULL.limbs(2);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_7dfc] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_7dfc_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_7dfc] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_7dfc_return_output := u320_t_NULL.limbs(0);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_7dfc] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_7dfc_return_output := u320_t_NULL.limbs(4);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_7dfc] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_7dfc_return_output := u320_t_NULL.limbs(1);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_7dfc_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_7dfc_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_7dfc_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_7dfc_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_7dfc_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_7a4b]_DUPLICATE_869a LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output := VAR_a.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_7a4b]_DUPLICATE_e228 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output := VAR_a.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_e477]_DUPLICATE_e531 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_e477]_DUPLICATE_226e LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_e477_DUPLICATE_226e_return_output := VAR_b.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_e477]_DUPLICATE_632a LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_e477_DUPLICATE_632a_return_output := VAR_b.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_7a4b]_DUPLICATE_5233 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_5233_return_output := VAR_a.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_7a4b]_DUPLICATE_acaf LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_acaf_return_output := VAR_a.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_e477]_DUPLICATE_2c13 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output := VAR_b.limbs(0);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_e477] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_e477_return_output := VAR_b.limbs(4);

     -- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_7a4b] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_7a4b_return_output := VAR_a.limbs(4);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_869a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_e477_DUPLICATE_2c13_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_e228_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_e477_DUPLICATE_e531_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_acaf_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_acaf_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_acaf_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_e477_DUPLICATE_632a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_e477_DUPLICATE_632a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_e477_DUPLICATE_632a_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_5233_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_7a4b_DUPLICATE_5233_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_e477_DUPLICATE_226e_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_e477_DUPLICATE_226e_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_e477_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_7a4b_return_output;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_7204] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_7204_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_product_poly1305_h_l127_c22_37c3_0;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_product_poly1305_h_l127_c22_37c3_0;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_2a7e] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_right;

     -- Write to comb signals
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_2a7e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l132_c21_fd3f_return_output;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8597] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8597_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_fec3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_fe6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_fe6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_09f7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_09f7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4c9a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_0a85] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_0a85_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_9973] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_9973_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_b459] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_b459_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_d7df] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_83f1] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_0285] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_right;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;

     -- Write to comb signals
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left := REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_0285_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_83f1_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_de17] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output;

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_de17_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_475c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_958d] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_42fd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_42fd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_866a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_ee02] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_ee02_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_866a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_1838] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_1838_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_5dcb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_0a27] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_0a27_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l131_c13_477c;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_5e22] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_9e29] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l132_c21_fd3f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_9e29_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_5e22_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l132_c21_fd3f_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_high_poly1305_h_l134_c13_c87d;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_3e3b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX[poly1305_h_l134_c22_c68b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_cond;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iftrue;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_3e3b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_MUX_poly1305_h_l134_c22_c68b_return_output;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_33f6] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_33f6_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_high_poly1305_h_l134_c13_c87d;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_886b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_886b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_low_poly1305_h_l133_c13_fd24;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_39a3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left := VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l131_c13_477c;
     -- FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_c44d] LATENCY=1
     -- Inputs
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_left;
     FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_right;

     -- Write to comb signals
     COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     -- Submodule outputs
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output := FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output;

     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 := resize(VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c44d_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_123a] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_123a_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24,
     VAR_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_123a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_fec3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4c9a_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_d7df_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE0_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     -- Stage 1
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_475c_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_958d_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_5dcb_right;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     REG_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left <= COMB_STAGE1_FOR_poly1305_h_l120_c5_47f7_ITER_4_FOR_poly1305_h_l123_c9_9e16_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_39a3_left;
     -- Stage 2
     REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_0_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_1_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_2_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
     REG_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24 <= COMB_STAGE2_FOR_poly1305_h_l120_c5_47f7_ITER_3_FOR_poly1305_h_l123_c9_9e16_ITER_0_low_poly1305_h_l133_c13_fd24;
 end if;
end process;

end arch;
