-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 16
entity axis128_keep_count_0CLK_08de2a73 is
port(
 axis : in axis128_t;
 return_output : out unsigned(4 downto 0));
end axis128_keep_count_0CLK_08de2a73;
architecture arch of axis128_keep_count_0CLK_08de2a73 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_72ee]
signal FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_bd78]
signal FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_dda2]
signal FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_541b]
signal FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_61e7]
signal FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_487b]
signal FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_b012]
signal FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_f642]
signal FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_c852]
signal FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_9625]
signal FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_9ef9]
signal FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_14a2]
signal FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_5364]
signal FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_dec9]
signal FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_d25f]
signal FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_0f08]
signal FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output : unsigned(5 downto 0);


begin

-- SUBMODULE INSTANCES 
-- FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left,
FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right,
FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left,
FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right,
FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left,
FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right,
FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left,
FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right,
FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left,
FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right,
FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left,
FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right,
FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left,
FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right,
FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left,
FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right,
FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left,
FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right,
FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left,
FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right,
FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left,
FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right,
FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left,
FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right,
FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left,
FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right,
FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left,
FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right,
FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left,
FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right,
FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output);

-- FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08 : 0 clocks latency
FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left,
FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right,
FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 axis,
 -- All submodule outputs
 FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output,
 FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(4 downto 0);
 variable VAR_axis : axis128_t;
 variable VAR_rv : unsigned(4 downto 0);
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_rv_axis_h_l91_c5_e15d : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_38c6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output : unsigned(5 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left := to_unsigned(0, 5);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_axis := axis;

     -- Submodule level 0
     -- FOR_axis_h_l90_c3_7bdd_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(11);

     -- FOR_axis_h_l90_c3_7bdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(0);

     -- FOR_axis_h_l90_c3_7bdd_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(6);

     -- FOR_axis_h_l90_c3_7bdd_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(8);

     -- FOR_axis_h_l90_c3_7bdd_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(3);

     -- FOR_axis_h_l90_c3_7bdd_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(9);

     -- FOR_axis_h_l90_c3_7bdd_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(13);

     -- FOR_axis_h_l90_c3_7bdd_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(10);

     -- FOR_axis_h_l90_c3_7bdd_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(7);

     -- FOR_axis_h_l90_c3_7bdd_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(14);

     -- FOR_axis_h_l90_c3_7bdd_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(5);

     -- FOR_axis_h_l90_c3_7bdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(2);

     -- FOR_axis_h_l90_c3_7bdd_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(12);

     -- FOR_axis_h_l90_c3_7bdd_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(4);

     -- FOR_axis_h_l90_c3_7bdd_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(15);

     -- FOR_axis_h_l90_c3_7bdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d[axis_h_l91_c11_38c6] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_38c6_return_output := VAR_axis.tkeep(1);

     -- Submodule level 1
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_38c6_return_output;
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right := VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_38c6_return_output;
     -- FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_72ee] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_left;
     FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output := FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output;

     -- Submodule level 2
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_72ee_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_0_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_bd78] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_left;
     FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output := FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output;

     -- Submodule level 3
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_bd78_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_1_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_dda2] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_left;
     FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output := FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output;

     -- Submodule level 4
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_dda2_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_2_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_541b] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_left;
     FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output := FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output;

     -- Submodule level 5
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_541b_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_3_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_61e7] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_left;
     FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output := FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output;

     -- Submodule level 6
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_61e7_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_4_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_487b] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_left;
     FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output := FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output;

     -- Submodule level 7
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_487b_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_5_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_b012] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_left;
     FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output := FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output;

     -- Submodule level 8
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_b012_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_6_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_f642] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_left;
     FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output := FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output;

     -- Submodule level 9
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_f642_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_7_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_c852] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_left;
     FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output := FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output;

     -- Submodule level 10
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_c852_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_8_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_9625] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_left;
     FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output := FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output;

     -- Submodule level 11
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_9625_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_9_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_9ef9] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_left;
     FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output := FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output;

     -- Submodule level 12
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_9ef9_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_10_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_14a2] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_left;
     FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output := FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output;

     -- Submodule level 13
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_14a2_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_11_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_5364] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_left;
     FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output := FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output;

     -- Submodule level 14
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_5364_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_12_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_dec9] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_left;
     FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output := FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output;

     -- Submodule level 15
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_dec9_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_13_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_d25f] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_left;
     FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output := FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output;

     -- Submodule level 16
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_d25f_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left := VAR_FOR_axis_h_l90_c3_7bdd_ITER_14_rv_axis_h_l91_c5_e15d;
     -- FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_0f08] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_left;
     FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right <= VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output := FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output;

     -- Submodule level 17
     VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_rv_axis_h_l91_c5_e15d := resize(VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_0f08_return_output, 5);
     VAR_return_output := VAR_FOR_axis_h_l90_c3_7bdd_ITER_15_rv_axis_h_l91_c5_e15d;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
