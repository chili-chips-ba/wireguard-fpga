-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.038461538461538464, 0.07692307692307693, 0.11538461538461539, 0.15384615384615385, 0.19230769230769232, 0.23076923076923078, 0.2692307692307693, 0.3076923076923077, 0.34615384615384615, 0.3846153846153846, 0.423076923076923, 0.46153846153846145, 0.4999999999999999, 0.5384615384615383, 0.5769230769230768, 0.6153846153846152, 0.6538461538461536, 0.6923076923076921, 0.7307692307692305, 0.7692307692307689, 0.8076923076923074, 0.8461538461538458, 0.8846153846153842, 0.9230769230769227, 0.9615384615384611]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 27
entity chacha20_block_25CLK_be909a13 is
port(
 clk : in std_logic;
 state : in chacha20_state;
 return_output : out chacha20_state);
end chacha20_block_25CLK_be909a13;
architecture arch of chacha20_block_25CLK_be909a13 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 25;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 1
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 2
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 3
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 4
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 5
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 6
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 7
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 8
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 9
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 10
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 11
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 12
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 13
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 14
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 15
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 16
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 17
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 18
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 19
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 20
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 21
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 22
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 23
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Stage 24
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
-- Each function instance gets signals
-- chacha20_block_step[chacha20_h_l72_c28_c4e8]
signal chacha20_block_step_chacha20_h_l72_c28_c4e8_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l73_c28_9045]
signal chacha20_block_step_chacha20_h_l73_c28_9045_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l73_c28_9045_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l74_c28_a3d4]
signal chacha20_block_step_chacha20_h_l74_c28_a3d4_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l75_c28_aab9]
signal chacha20_block_step_chacha20_h_l75_c28_aab9_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l75_c28_aab9_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l76_c28_fed3]
signal chacha20_block_step_chacha20_h_l76_c28_fed3_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l76_c28_fed3_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l77_c28_ecce]
signal chacha20_block_step_chacha20_h_l77_c28_ecce_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l77_c28_ecce_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l78_c28_25fc]
signal chacha20_block_step_chacha20_h_l78_c28_25fc_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l78_c28_25fc_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l79_c28_ffaf]
signal chacha20_block_step_chacha20_h_l79_c28_ffaf_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l80_c28_6d70]
signal chacha20_block_step_chacha20_h_l80_c28_6d70_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l80_c28_6d70_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l81_c29_5148]
signal chacha20_block_step_chacha20_h_l81_c29_5148_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l81_c29_5148_return_output : chacha20_state;

-- FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_b94b]
signal FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);

function CONST_REF_RD_chacha20_state_chacha20_state_23da( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return chacha20_state is
 
  variable base : chacha20_state; 
  variable return_output : chacha20_state;
begin
      base.state(0) := ref_toks_0;
      base.state(1) := ref_toks_1;
      base.state(2) := ref_toks_2;
      base.state(3) := ref_toks_3;
      base.state(4) := ref_toks_4;
      base.state(5) := ref_toks_5;
      base.state(6) := ref_toks_6;
      base.state(7) := ref_toks_7;
      base.state(8) := ref_toks_8;
      base.state(9) := ref_toks_9;
      base.state(10) := ref_toks_10;
      base.state(11) := ref_toks_11;
      base.state(12) := ref_toks_12;
      base.state(13) := ref_toks_13;
      base.state(14) := ref_toks_14;
      base.state(15) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- chacha20_block_step_chacha20_h_l72_c28_c4e8 : 2 clocks latency
chacha20_block_step_chacha20_h_l72_c28_c4e8 : entity work.chacha20_block_step_2CLK_9dedafab port map (
clk,
chacha20_block_step_chacha20_h_l72_c28_c4e8_state0,
chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output);

-- chacha20_block_step_chacha20_h_l73_c28_9045 : 3 clocks latency
chacha20_block_step_chacha20_h_l73_c28_9045 : entity work.chacha20_block_step_3CLK_0846ca6c port map (
clk,
chacha20_block_step_chacha20_h_l73_c28_9045_state0,
chacha20_block_step_chacha20_h_l73_c28_9045_return_output);

-- chacha20_block_step_chacha20_h_l74_c28_a3d4 : 2 clocks latency
chacha20_block_step_chacha20_h_l74_c28_a3d4 : entity work.chacha20_block_step_2CLK_a128b32a port map (
clk,
chacha20_block_step_chacha20_h_l74_c28_a3d4_state0,
chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output);

-- chacha20_block_step_chacha20_h_l75_c28_aab9 : 3 clocks latency
chacha20_block_step_chacha20_h_l75_c28_aab9 : entity work.chacha20_block_step_3CLK_b0a08188 port map (
clk,
chacha20_block_step_chacha20_h_l75_c28_aab9_state0,
chacha20_block_step_chacha20_h_l75_c28_aab9_return_output);

-- chacha20_block_step_chacha20_h_l76_c28_fed3 : 2 clocks latency
chacha20_block_step_chacha20_h_l76_c28_fed3 : entity work.chacha20_block_step_2CLK_b472b82d port map (
clk,
chacha20_block_step_chacha20_h_l76_c28_fed3_state0,
chacha20_block_step_chacha20_h_l76_c28_fed3_return_output);

-- chacha20_block_step_chacha20_h_l77_c28_ecce : 3 clocks latency
chacha20_block_step_chacha20_h_l77_c28_ecce : entity work.chacha20_block_step_3CLK_9b7a5add port map (
clk,
chacha20_block_step_chacha20_h_l77_c28_ecce_state0,
chacha20_block_step_chacha20_h_l77_c28_ecce_return_output);

-- chacha20_block_step_chacha20_h_l78_c28_25fc : 2 clocks latency
chacha20_block_step_chacha20_h_l78_c28_25fc : entity work.chacha20_block_step_2CLK_b6cd9d54 port map (
clk,
chacha20_block_step_chacha20_h_l78_c28_25fc_state0,
chacha20_block_step_chacha20_h_l78_c28_25fc_return_output);

-- chacha20_block_step_chacha20_h_l79_c28_ffaf : 3 clocks latency
chacha20_block_step_chacha20_h_l79_c28_ffaf : entity work.chacha20_block_step_3CLK_7f7fdb6d port map (
clk,
chacha20_block_step_chacha20_h_l79_c28_ffaf_state0,
chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output);

-- chacha20_block_step_chacha20_h_l80_c28_6d70 : 3 clocks latency
chacha20_block_step_chacha20_h_l80_c28_6d70 : entity work.chacha20_block_step_3CLK_d12c72c2 port map (
clk,
chacha20_block_step_chacha20_h_l80_c28_6d70_state0,
chacha20_block_step_chacha20_h_l80_c28_6d70_return_output);

-- chacha20_block_step_chacha20_h_l81_c29_5148 : 2 clocks latency
chacha20_block_step_chacha20_h_l81_c29_5148 : entity work.chacha20_block_step_2CLK_a1536939 port map (
clk,
chacha20_block_step_chacha20_h_l81_c29_5148_state0,
chacha20_block_step_chacha20_h_l81_c29_5148_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);

-- FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : 0 clocks latency
FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left,
FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 state,
 -- Registers
 -- Stage 0
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 1
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 2
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 3
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 4
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 5
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 6
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 7
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 8
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 9
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 10
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 11
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 12
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 13
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 14
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 15
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 16
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 17
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 18
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 19
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 20
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 21
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 22
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 23
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- Stage 24
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right,
 -- All submodule outputs
 chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output,
 chacha20_block_step_chacha20_h_l73_c28_9045_return_output,
 chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output,
 chacha20_block_step_chacha20_h_l75_c28_aab9_return_output,
 chacha20_block_step_chacha20_h_l76_c28_fed3_return_output,
 chacha20_block_step_chacha20_h_l77_c28_ecce_return_output,
 chacha20_block_step_chacha20_h_l78_c28_25fc_return_output,
 chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output,
 chacha20_block_step_chacha20_h_l80_c28_6d70_return_output,
 chacha20_block_step_chacha20_h_l81_c29_5148_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output,
 FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : chacha20_state;
 variable VAR_state : chacha20_state;
 variable VAR_output : chacha20_state;
 variable VAR_step1 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output : chacha20_state;
 variable VAR_step2 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_9045_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_9045_return_output : chacha20_state;
 variable VAR_step3 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output : chacha20_state;
 variable VAR_step4 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_return_output : chacha20_state;
 variable VAR_step5 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_return_output : chacha20_state;
 variable VAR_step6 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_return_output : chacha20_state;
 variable VAR_step7 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_return_output : chacha20_state;
 variable VAR_step8 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output : chacha20_state;
 variable VAR_step9 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_return_output : chacha20_state;
 variable VAR_step10 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_5148_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output : chacha20_state;
 variable VAR_i : unsigned(3 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_output_state_0_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_output_state_1_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_output_state_2_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_output_state_3_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_output_state_4_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_output_state_5_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_output_state_6_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_output_state_7_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_output_state_8_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_output_state_9_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_output_state_10_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_output_state_11_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_output_state_12_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_output_state_13_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_output_state_14_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_output_state_15_chacha20_h_l87_c9_0fc6 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_9098_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f9af_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_870e_return_output : chacha20_state;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_state := state;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_state0 := VAR_state;
     -- FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(7);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(9);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(14);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(2);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(6);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(0);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(3);

     -- chacha20_block_step[chacha20_h_l72_c28_c4e8] LATENCY=2
     -- Inputs
     chacha20_block_step_chacha20_h_l72_c28_c4e8_state0 <= VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_state0;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(13);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(12);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(10);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(1);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(15);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(5);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(8);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(4);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c45_f9af] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f9af_return_output := VAR_state.state(11);

     -- Submodule level 1
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_f9af_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_f9af_return_output;
     -- Write to comb signals
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output := chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l73_c28_9045_state0 := VAR_chacha20_block_step_chacha20_h_l72_c28_c4e8_return_output;
     -- chacha20_block_step[chacha20_h_l73_c28_9045] LATENCY=3
     -- Inputs
     chacha20_block_step_chacha20_h_l73_c28_9045_state0 <= VAR_chacha20_block_step_chacha20_h_l73_c28_9045_state0;

     -- Write to comb signals
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l73_c28_9045_return_output := chacha20_block_step_chacha20_h_l73_c28_9045_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_state0 := VAR_chacha20_block_step_chacha20_h_l73_c28_9045_return_output;
     -- chacha20_block_step[chacha20_h_l74_c28_a3d4] LATENCY=2
     -- Inputs
     chacha20_block_step_chacha20_h_l74_c28_a3d4_state0 <= VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_state0;

     -- Write to comb signals
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output := chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_state0 := VAR_chacha20_block_step_chacha20_h_l74_c28_a3d4_return_output;
     -- chacha20_block_step[chacha20_h_l75_c28_aab9] LATENCY=3
     -- Inputs
     chacha20_block_step_chacha20_h_l75_c28_aab9_state0 <= VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_state0;

     -- Write to comb signals
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_return_output := chacha20_block_step_chacha20_h_l75_c28_aab9_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_state0 := VAR_chacha20_block_step_chacha20_h_l75_c28_aab9_return_output;
     -- chacha20_block_step[chacha20_h_l76_c28_fed3] LATENCY=2
     -- Inputs
     chacha20_block_step_chacha20_h_l76_c28_fed3_state0 <= VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_state0;

     -- Write to comb signals
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_return_output := chacha20_block_step_chacha20_h_l76_c28_fed3_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_state0 := VAR_chacha20_block_step_chacha20_h_l76_c28_fed3_return_output;
     -- chacha20_block_step[chacha20_h_l77_c28_ecce] LATENCY=3
     -- Inputs
     chacha20_block_step_chacha20_h_l77_c28_ecce_state0 <= VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_state0;

     -- Write to comb signals
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_return_output := chacha20_block_step_chacha20_h_l77_c28_ecce_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_state0 := VAR_chacha20_block_step_chacha20_h_l77_c28_ecce_return_output;
     -- chacha20_block_step[chacha20_h_l78_c28_25fc] LATENCY=2
     -- Inputs
     chacha20_block_step_chacha20_h_l78_c28_25fc_state0 <= VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_state0;

     -- Write to comb signals
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_return_output := chacha20_block_step_chacha20_h_l78_c28_25fc_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_state0 := VAR_chacha20_block_step_chacha20_h_l78_c28_25fc_return_output;
     -- chacha20_block_step[chacha20_h_l79_c28_ffaf] LATENCY=3
     -- Inputs
     chacha20_block_step_chacha20_h_l79_c28_ffaf_state0 <= VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_state0;

     -- Write to comb signals
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output := chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_state0 := VAR_chacha20_block_step_chacha20_h_l79_c28_ffaf_return_output;
     -- chacha20_block_step[chacha20_h_l80_c28_6d70] LATENCY=3
     -- Inputs
     chacha20_block_step_chacha20_h_l80_c28_6d70_state0 <= VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_state0;

     -- Write to comb signals
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_return_output := chacha20_block_step_chacha20_h_l80_c28_6d70_return_output;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l81_c29_5148_state0 := VAR_chacha20_block_step_chacha20_h_l80_c28_6d70_return_output;
     -- chacha20_block_step[chacha20_h_l81_c29_5148] LATENCY=2
     -- Inputs
     chacha20_block_step_chacha20_h_l81_c29_5148_state0 <= VAR_chacha20_block_step_chacha20_h_l81_c29_5148_state0;

     -- Write to comb signals
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;

     -- Write to comb signals
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right := REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Submodule outputs
     VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output := chacha20_block_step_chacha20_h_l81_c29_5148_return_output;

     -- Submodule level 0
     -- FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(3);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(11);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(5);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(0);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(4);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(12);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(9);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(14);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(7);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(8);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(1);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(2);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(13);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(15);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(6);

     -- FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c27_9098] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_9098_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_5148_return_output.state(10);

     -- Submodule level 1
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_9098_return_output;
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left := VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_9098_return_output;
     -- FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_b94b] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_left;
     FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output := FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output;

     -- Submodule level 2
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_output_state_0_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_output_state_10_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_output_state_11_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_output_state_12_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_output_state_13_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_output_state_14_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_output_state_15_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_output_state_1_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_output_state_2_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_output_state_3_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_output_state_4_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_output_state_5_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_output_state_6_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_output_state_7_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_output_state_8_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_output_state_9_chacha20_h_l87_c9_0fc6 := resize(VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_return_output, 32);
     -- CONST_REF_RD_chacha20_state_chacha20_state_23da[chacha20_h_l90_c12_870e] LATENCY=0
     VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_870e_return_output := CONST_REF_RD_chacha20_state_chacha20_state_23da(
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_0_output_state_0_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_1_output_state_1_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_2_output_state_2_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_3_output_state_3_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_4_output_state_4_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_5_output_state_5_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_6_output_state_6_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_7_output_state_7_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_8_output_state_8_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_9_output_state_9_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_10_output_state_10_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_11_output_state_11_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_12_output_state_12_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_13_output_state_13_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_14_output_state_14_chacha20_h_l87_c9_0fc6,
     VAR_FOR_chacha20_h_l85_c5_25c4_ITER_15_output_state_15_chacha20_h_l87_c9_0fc6);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_870e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE0_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 1
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE1_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 2
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE2_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 3
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE3_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 4
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE4_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 5
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE5_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 6
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE6_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 7
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE7_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 8
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE8_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 9
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE9_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 10
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE10_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 11
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE11_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 12
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE12_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 13
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE13_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 14
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE14_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 15
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE15_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 16
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE16_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 17
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE17_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 18
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE18_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 19
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE19_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 20
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE20_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 21
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE21_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 22
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE22_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 23
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE23_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     -- Stage 24
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
     REG_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right <= COMB_STAGE24_FOR_chacha20_h_l85_c5_25c4_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_b94b_right;
 end if;
end process;

end arch;
