mem['h0000] = 32'h00000517;
mem['h0001] = 32'h7A850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h60C18593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h2A0000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'h6081A703;
mem['h001D] = 32'h100007B7;
mem['h001E] = 32'h60878793;
mem['h001F] = 32'h00F707B3;
mem['h0020] = 32'h00A70733;
mem['h0021] = 32'h60E1A423;
mem['h0022] = 32'h000016B7;
mem['h0023] = 32'h80068693;
mem['h0024] = 32'h00E6D463;
mem['h0025] = 32'h00100073;
mem['h0026] = 32'h00078513;
mem['h0027] = 32'h00008067;
mem['h0028] = 32'h00052783;
mem['h0029] = 32'h0007A783;
mem['h002A] = 32'h0187A783;
mem['h002B] = 32'h0007A783;
mem['h002C] = 32'h0007A783;
mem['h002D] = 32'h0017F793;
mem['h002E] = 32'h20078463;
mem['h002F] = 32'h00052783;
mem['h0030] = 32'h100006B7;
mem['h0031] = 32'h00068613;
mem['h0032] = 32'h0007A783;
mem['h0033] = 32'h00064703;
mem['h0034] = 32'hFFFF08B7;
mem['h0035] = 32'h0107A783;
mem['h0036] = 32'h00777713;
mem['h0037] = 32'h0007A583;
mem['h0038] = 32'h0005A783;
mem['h0039] = 32'hFF87F793;
mem['h003A] = 32'h00E7E7B3;
mem['h003B] = 32'h00F5A023;
mem['h003C] = 32'h00052783;
mem['h003D] = 32'h00164703;
mem['h003E] = 32'h0007A783;
mem['h003F] = 32'h00777713;
mem['h0040] = 32'h00371713;
mem['h0041] = 32'h0107A783;
mem['h0042] = 32'h0007A583;
mem['h0043] = 32'h0005A783;
mem['h0044] = 32'hFC77F793;
mem['h0045] = 32'h00E7E7B3;
mem['h0046] = 32'h00F5A023;
mem['h0047] = 32'h00052783;
mem['h0048] = 32'h00264703;
mem['h0049] = 32'h0007A783;
mem['h004A] = 32'h00177713;
mem['h004B] = 32'h00671713;
mem['h004C] = 32'h0107A783;
mem['h004D] = 32'h0007A583;
mem['h004E] = 32'h0005A783;
mem['h004F] = 32'hFBF7F793;
mem['h0050] = 32'h00E7E7B3;
mem['h0051] = 32'h00F5A023;
mem['h0052] = 32'h00052783;
mem['h0053] = 32'h00364703;
mem['h0054] = 32'h0007A783;
mem['h0055] = 32'h00177713;
mem['h0056] = 32'h00771713;
mem['h0057] = 32'h0107A783;
mem['h0058] = 32'h0007A583;
mem['h0059] = 32'h0005A783;
mem['h005A] = 32'hF7F7F793;
mem['h005B] = 32'h00E7E7B3;
mem['h005C] = 32'h00F5A023;
mem['h005D] = 32'hFFFF85B7;
mem['h005E] = 32'h00068713;
mem['h005F] = 32'h00000793;
mem['h0060] = 32'h00068693;
mem['h0061] = 32'hFFF58593;
mem['h0062] = 32'h00052603;
mem['h0063] = 32'h00872803;
mem['h0064] = 32'h01078793;
mem['h0065] = 32'h00062603;
mem['h0066] = 32'h01070713;
mem['h0067] = 32'h00062603;
mem['h0068] = 32'h00062603;
mem['h0069] = 32'h01062023;
mem['h006A] = 32'h00052603;
mem['h006B] = 32'hFFC72803;
mem['h006C] = 32'h00062603;
mem['h006D] = 32'h00462603;
mem['h006E] = 32'h00062603;
mem['h006F] = 32'h01062023;
mem['h0070] = 32'h00052603;
mem['h0071] = 32'h00072803;
mem['h0072] = 32'h00062603;
mem['h0073] = 32'h00862603;
mem['h0074] = 32'h00062603;
mem['h0075] = 32'h01062023;
mem['h0076] = 32'h00052603;
mem['h0077] = 32'h00472803;
mem['h0078] = 32'h00062603;
mem['h0079] = 32'h00C62603;
mem['h007A] = 32'h00062603;
mem['h007B] = 32'h01062023;
mem['h007C] = 32'h0046A803;
mem['h007D] = 32'h0507FE63;
mem['h007E] = 32'h00052603;
mem['h007F] = 32'h00062603;
mem['h0080] = 32'h01062603;
mem['h0081] = 32'h00062803;
mem['h0082] = 32'h00082603;
mem['h0083] = 32'h01166633;
mem['h0084] = 32'h00C82023;
mem['h0085] = 32'h00052603;
mem['h0086] = 32'h00062603;
mem['h0087] = 32'h01062603;
mem['h0088] = 32'h00062803;
mem['h0089] = 32'h00082603;
mem['h008A] = 32'h00B67633;
mem['h008B] = 32'h00C82023;
mem['h008C] = 32'h00052603;
mem['h008D] = 32'h00062603;
mem['h008E] = 32'h01462603;
mem['h008F] = 32'h00062803;
mem['h0090] = 32'h00082603;
mem['h0091] = 32'h00166613;
mem['h0092] = 32'h00C82023;
mem['h0093] = 32'hF3DFF06F;
mem['h0094] = 32'h00052703;
mem['h0095] = 32'h000106B7;
mem['h0096] = 32'hFFF68693;
mem['h0097] = 32'h00072703;
mem['h0098] = 32'h410787B3;
mem['h0099] = 32'h40F6D7B3;
mem['h009A] = 32'h01072703;
mem['h009B] = 32'h01079793;
mem['h009C] = 32'h00072603;
mem['h009D] = 32'h00062703;
mem['h009E] = 32'h00D77733;
mem['h009F] = 32'h00F767B3;
mem['h00A0] = 32'h00F62023;
mem['h00A1] = 32'h00052783;
mem['h00A2] = 32'h000086B7;
mem['h00A3] = 32'h0007A783;
mem['h00A4] = 32'h0107A783;
mem['h00A5] = 32'h0007A703;
mem['h00A6] = 32'h00072783;
mem['h00A7] = 32'h00D7E7B3;
mem['h00A8] = 32'h00F72023;
mem['h00A9] = 32'h00052783;
mem['h00AA] = 32'h0007A783;
mem['h00AB] = 32'h0147A783;
mem['h00AC] = 32'h0007A703;
mem['h00AD] = 32'h00072783;
mem['h00AE] = 32'h0017E793;
mem['h00AF] = 32'h00F72023;
mem['h00B0] = 32'h00008067;
mem['h00B1] = 32'h0FF5F593;
mem['h00B2] = 32'h00000793;
mem['h00B3] = 32'h00C79463;
mem['h00B4] = 32'h00008067;
mem['h00B5] = 32'h00F50733;
mem['h00B6] = 32'h00B70023;
mem['h00B7] = 32'h00178793;
mem['h00B8] = 32'hFEDFF06F;
mem['h00B9] = 32'h00000793;
mem['h00BA] = 32'h00C79463;
mem['h00BB] = 32'h00008067;
mem['h00BC] = 32'h00F58733;
mem['h00BD] = 32'h00074683;
mem['h00BE] = 32'h00F50733;
mem['h00BF] = 32'h00178793;
mem['h00C0] = 32'h00D70023;
mem['h00C1] = 32'hFE5FF06F;
mem['h00C2] = 32'hFE010113;
mem['h00C3] = 32'h02800513;
mem['h00C4] = 32'h00112E23;
mem['h00C5] = 32'h00812C23;
mem['h00C6] = 32'h00912A23;
mem['h00C7] = 32'h01212823;
mem['h00C8] = 32'h01312623;
mem['h00C9] = 32'h01412423;
mem['h00CA] = 32'h01512223;
mem['h00CB] = 32'hD45FF0EF;
mem['h00CC] = 32'h00050413;
mem['h00CD] = 32'h00800513;
mem['h00CE] = 32'hD39FF0EF;
mem['h00CF] = 32'h00050913;
mem['h00D0] = 32'h01C00513;
mem['h00D1] = 32'hD2DFF0EF;
mem['h00D2] = 32'h00050493;
mem['h00D3] = 32'h00400513;
mem['h00D4] = 32'hD21FF0EF;
mem['h00D5] = 32'h200007B7;
mem['h00D6] = 32'h00F52023;
mem['h00D7] = 32'h00A4A023;
mem['h00D8] = 32'h00400513;
mem['h00D9] = 32'hD0DFF0EF;
mem['h00DA] = 32'h200007B7;
mem['h00DB] = 32'h00478793;
mem['h00DC] = 32'h00F52023;
mem['h00DD] = 32'h00A4A223;
mem['h00DE] = 32'h00400513;
mem['h00DF] = 32'hCF5FF0EF;
mem['h00E0] = 32'h200007B7;
mem['h00E1] = 32'h00878793;
mem['h00E2] = 32'h00F52023;
mem['h00E3] = 32'h00A4A423;
mem['h00E4] = 32'h00400513;
mem['h00E5] = 32'hCDDFF0EF;
mem['h00E6] = 32'h200007B7;
mem['h00E7] = 32'h00C78793;
mem['h00E8] = 32'h00F52023;
mem['h00E9] = 32'h00A4A623;
mem['h00EA] = 32'h00400513;
mem['h00EB] = 32'hCC5FF0EF;
mem['h00EC] = 32'h200007B7;
mem['h00ED] = 32'h01078793;
mem['h00EE] = 32'h00F52023;
mem['h00EF] = 32'h00A4A823;
mem['h00F0] = 32'h00400513;
mem['h00F1] = 32'hCADFF0EF;
mem['h00F2] = 32'h200007B7;
mem['h00F3] = 32'h01478793;
mem['h00F4] = 32'h00F52023;
mem['h00F5] = 32'h00A4AA23;
mem['h00F6] = 32'h00400513;
mem['h00F7] = 32'hC95FF0EF;
mem['h00F8] = 32'h200007B7;
mem['h00F9] = 32'h01878793;
mem['h00FA] = 32'h00F52023;
mem['h00FB] = 32'h00A4AC23;
mem['h00FC] = 32'h00992023;
mem['h00FD] = 32'h01C00513;
mem['h00FE] = 32'hC79FF0EF;
mem['h00FF] = 32'h00050493;
mem['h0100] = 32'h00400513;
mem['h0101] = 32'hC6DFF0EF;
mem['h0102] = 32'h200007B7;
mem['h0103] = 32'h01C78793;
mem['h0104] = 32'h00F52023;
mem['h0105] = 32'h00A4A023;
mem['h0106] = 32'h00400513;
mem['h0107] = 32'hC55FF0EF;
mem['h0108] = 32'h200007B7;
mem['h0109] = 32'h02078793;
mem['h010A] = 32'h00F52023;
mem['h010B] = 32'h00A4A223;
mem['h010C] = 32'h00400513;
mem['h010D] = 32'hC3DFF0EF;
mem['h010E] = 32'h200007B7;
mem['h010F] = 32'h02478793;
mem['h0110] = 32'h00F52023;
mem['h0111] = 32'h00A4A423;
mem['h0112] = 32'h00400513;
mem['h0113] = 32'hC25FF0EF;
mem['h0114] = 32'h200007B7;
mem['h0115] = 32'h02878793;
mem['h0116] = 32'h00F52023;
mem['h0117] = 32'h00A4A623;
mem['h0118] = 32'h00400513;
mem['h0119] = 32'hC0DFF0EF;
mem['h011A] = 32'h200007B7;
mem['h011B] = 32'h02C78793;
mem['h011C] = 32'h00F52023;
mem['h011D] = 32'h00A4A823;
mem['h011E] = 32'h00400513;
mem['h011F] = 32'hBF5FF0EF;
mem['h0120] = 32'h200007B7;
mem['h0121] = 32'h03078793;
mem['h0122] = 32'h00F52023;
mem['h0123] = 32'h00A4AA23;
mem['h0124] = 32'h00400513;
mem['h0125] = 32'hBDDFF0EF;
mem['h0126] = 32'h200007B7;
mem['h0127] = 32'h03478793;
mem['h0128] = 32'h00F52023;
mem['h0129] = 32'h00A4AC23;
mem['h012A] = 32'h00992223;
mem['h012B] = 32'h01242023;
mem['h012C] = 32'h01000513;
mem['h012D] = 32'hBBDFF0EF;
mem['h012E] = 32'h00050493;
mem['h012F] = 32'h00400513;
mem['h0130] = 32'hBB1FF0EF;
mem['h0131] = 32'h200007B7;
mem['h0132] = 32'h03878793;
mem['h0133] = 32'h00F52023;
mem['h0134] = 32'h00A4A023;
mem['h0135] = 32'h00400513;
mem['h0136] = 32'hB99FF0EF;
mem['h0137] = 32'h200007B7;
mem['h0138] = 32'h03C78793;
mem['h0139] = 32'h00F52023;
mem['h013A] = 32'h00A4A223;
mem['h013B] = 32'h00400513;
mem['h013C] = 32'hB81FF0EF;
mem['h013D] = 32'h200007B7;
mem['h013E] = 32'h04078793;
mem['h013F] = 32'h00F52023;
mem['h0140] = 32'h00A4A423;
mem['h0141] = 32'h00400513;
mem['h0142] = 32'hB69FF0EF;
mem['h0143] = 32'h200007B7;
mem['h0144] = 32'h04478793;
mem['h0145] = 32'h00F52023;
mem['h0146] = 32'h00A4A623;
mem['h0147] = 32'h00942223;
mem['h0148] = 32'h00400513;
mem['h0149] = 32'hB4DFF0EF;
mem['h014A] = 32'h200007B7;
mem['h014B] = 32'h04878793;
mem['h014C] = 32'h00F52023;
mem['h014D] = 32'h200004B7;
mem['h014E] = 32'h200009B7;
mem['h014F] = 32'h00A42423;
mem['h0150] = 32'h00C40A13;
mem['h0151] = 32'h04C48493;
mem['h0152] = 32'h07C98993;
mem['h0153] = 32'h00C00513;
mem['h0154] = 32'hB21FF0EF;
mem['h0155] = 32'h00050913;
mem['h0156] = 32'h00400513;
mem['h0157] = 32'hB15FF0EF;
mem['h0158] = 32'h00952023;
mem['h0159] = 32'h00A92023;
mem['h015A] = 32'h00400513;
mem['h015B] = 32'hB05FF0EF;
mem['h015C] = 32'h00448793;
mem['h015D] = 32'h00F52023;
mem['h015E] = 32'h00A92223;
mem['h015F] = 32'h00400513;
mem['h0160] = 32'hAF1FF0EF;
mem['h0161] = 32'h00848793;
mem['h0162] = 32'h00F52023;
mem['h0163] = 32'h00A92423;
mem['h0164] = 32'h012A2023;
mem['h0165] = 32'h00C48493;
mem['h0166] = 32'h004A0A13;
mem['h0167] = 32'hFB3498E3;
mem['h0168] = 32'h00400513;
mem['h0169] = 32'hACDFF0EF;
mem['h016A] = 32'h00050913;
mem['h016B] = 32'h00400513;
mem['h016C] = 32'hAC1FF0EF;
mem['h016D] = 32'h00952023;
mem['h016E] = 32'h00A92023;
mem['h016F] = 32'h01242E23;
mem['h0170] = 32'h00400513;
mem['h0171] = 32'hAADFF0EF;
mem['h0172] = 32'h200007B7;
mem['h0173] = 32'h08078793;
mem['h0174] = 32'h00F52023;
mem['h0175] = 32'h02A42023;
mem['h0176] = 32'h00400513;
mem['h0177] = 32'hA95FF0EF;
mem['h0178] = 32'h200007B7;
mem['h0179] = 32'h08478793;
mem['h017A] = 32'h00F52023;
mem['h017B] = 32'h100004B7;
mem['h017C] = 32'h02A42223;
mem['h017D] = 32'h00048493;
mem['h017E] = 32'h5F000993;
mem['h017F] = 32'h60000A13;
mem['h0180] = 32'h00100A93;
mem['h0181] = 32'h00200913;
mem['h0182] = 32'h00048023;
mem['h0183] = 32'h00049123;
mem['h0184] = 32'h00042783;
mem['h0185] = 32'h0047A783;
mem['h0186] = 32'h0187A783;
mem['h0187] = 32'h0007A783;
mem['h0188] = 32'h0007A783;
mem['h0189] = 32'h0017F793;
mem['h018A] = 32'h0E078E63;
mem['h018B] = 32'h00042783;
mem['h018C] = 32'h00048713;
mem['h018D] = 32'h0047A783;
mem['h018E] = 32'h0107A783;
mem['h018F] = 32'h0007A783;
mem['h0190] = 32'h0007A783;
mem['h0191] = 32'h0037D793;
mem['h0192] = 32'h0077F793;
mem['h0193] = 32'h00F480A3;
mem['h0194] = 32'h00000793;
mem['h0195] = 32'h06F9E263;
mem['h0196] = 32'h00042683;
mem['h0197] = 32'h0046A683;
mem['h0198] = 32'h0006A683;
mem['h0199] = 32'h0006A683;
mem['h019A] = 32'h0006A683;
mem['h019B] = 32'h00D72423;
mem['h019C] = 32'h00042683;
mem['h019D] = 32'h0046A683;
mem['h019E] = 32'h0046A683;
mem['h019F] = 32'h0006A683;
mem['h01A0] = 32'h0006A683;
mem['h01A1] = 32'h00D72623;
mem['h01A2] = 32'h00042683;
mem['h01A3] = 32'h0046A683;
mem['h01A4] = 32'h0086A683;
mem['h01A5] = 32'h0006A683;
mem['h01A6] = 32'h0006A683;
mem['h01A7] = 32'h00D72823;
mem['h01A8] = 32'h00042683;
mem['h01A9] = 32'h0046A683;
mem['h01AA] = 32'h00C6A683;
mem['h01AB] = 32'h0006A683;
mem['h01AC] = 32'h0006A683;
mem['h01AD] = 32'h00D72A23;
mem['h01AE] = 32'h00042683;
mem['h01AF] = 32'h01070713;
mem['h01B0] = 32'h0046A683;
mem['h01B1] = 32'h0106A683;
mem['h01B2] = 32'h0006A683;
mem['h01B3] = 32'h0006A683;
mem['h01B4] = 32'h01069613;
mem['h01B5] = 32'h06065A63;
mem['h01B6] = 32'h00042703;
mem['h01B7] = 32'h00472703;
mem['h01B8] = 32'h01072703;
mem['h01B9] = 32'h00072703;
mem['h01BA] = 32'h00275703;
mem['h01BB] = 32'h00177693;
mem['h01BC] = 32'h04069663;
mem['h01BD] = 32'h00FA7463;
mem['h01BE] = 32'h60000793;
mem['h01BF] = 32'h00F4A223;
mem['h01C0] = 32'h00042783;
mem['h01C1] = 32'h0047A783;
mem['h01C2] = 32'h0147A783;
mem['h01C3] = 32'h0007A703;
mem['h01C4] = 32'h00072783;
mem['h01C5] = 32'h0017E793;
mem['h01C6] = 32'h00F72023;
mem['h01C7] = 32'h0044A783;
mem['h01C8] = 32'h04079663;
mem['h01C9] = 32'h00842783;
mem['h01CA] = 32'h0007A703;
mem['h01CB] = 32'h00072783;
mem['h01CC] = 32'hDFF7F793;
mem['h01CD] = 32'h00F72023;
mem['h01CE] = 32'hED1FF06F;
mem['h01CF] = 32'h00178793;
mem['h01D0] = 32'h00175713;
mem['h01D1] = 32'hFA9FF06F;
mem['h01D2] = 32'h00042683;
mem['h01D3] = 32'h01078793;
mem['h01D4] = 32'h0046A683;
mem['h01D5] = 32'h0146A683;
mem['h01D6] = 32'h0006A603;
mem['h01D7] = 32'h00062683;
mem['h01D8] = 32'h0016E693;
mem['h01D9] = 32'h00D62023;
mem['h01DA] = 32'hEEDFF06F;
mem['h01DB] = 32'h00842783;
mem['h01DC] = 32'h0007A703;
mem['h01DD] = 32'h00072783;
mem['h01DE] = 32'h2007E793;
mem['h01DF] = 32'h00F72023;
mem['h01E0] = 32'h0014C783;
mem['h01E1] = 32'h01579C63;
mem['h01E2] = 32'h01248023;
mem['h01E3] = 32'h00040513;
mem['h01E4] = 32'h015481A3;
mem['h01E5] = 32'h90DFF0EF;
mem['h01E6] = 32'hE71FF06F;
mem['h01E7] = 32'hE72796E3;
mem['h01E8] = 32'h01548023;
mem['h01E9] = 32'hFE9FF06F;
