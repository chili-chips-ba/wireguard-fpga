-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_0CLK_babc4282 is
port(
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_0CLK_babc4282;
architecture arch of uint320_mul_0CLK_babc4282 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_27b4]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_e7fe]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6486]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_8f00]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4669]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_001b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_302c]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_8e84]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_c4ed]
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_61d2]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8e6c]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6eed]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_c84f]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_b299]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_6a38]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_fc1c]
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d7f4]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_683c]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_42ab]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_4553]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_a9da]
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_91bb]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_d037]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6e6c]
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a]
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7]
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_38af]
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right,
FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right,
FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right,
FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5 : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right,
FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output);

-- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af : 0 clocks latency
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right,
FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output,
 FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_df2e_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_df2e_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_df2e_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_df2e_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3d65_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_df2e_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_93a3_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_3224_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_35b8_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6eb6_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_610e_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_3684_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse := to_unsigned(0, 64);
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_df2e] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_df2e_return_output := u320_t_NULL.limbs(0);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_df2e] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_df2e_return_output := u320_t_NULL.limbs(2);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_df2e] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_df2e_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_df2e] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_df2e_return_output := u320_t_NULL.limbs(4);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_df2e] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_df2e_return_output := u320_t_NULL.limbs(1);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_df2e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_df2e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_df2e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_df2e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_df2e_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_93a3]_DUPLICATE_610e LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_610e_return_output := VAR_a.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_93a3]_DUPLICATE_478a LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output := VAR_a.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_93a3]_DUPLICATE_89ce LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output := VAR_a.limbs(0);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_93a3] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_93a3_return_output := VAR_a.limbs(4);

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_3d65] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3d65_return_output := VAR_b.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_3d65]_DUPLICATE_35b8 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_35b8_return_output := VAR_b.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_3d65]_DUPLICATE_6c74 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output := VAR_b.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_3d65]_DUPLICATE_00c7 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_93a3]_DUPLICATE_3684 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_3684_return_output := VAR_a.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_3d65]_DUPLICATE_6eb6 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6eb6_return_output := VAR_b.limbs(3);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_89ce_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6c74_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_478a_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_00c7_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_610e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_610e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_610e_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_35b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_35b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_35b8_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_3684_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_93a3_DUPLICATE_3684_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6eb6_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_3d65_DUPLICATE_6eb6_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_3d65_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_93a3_return_output;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_0f6a] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_0f6a_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_product_poly1305_h_l127_c22_85bf_0;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_product_poly1305_h_l127_c22_85bf_0;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_27b4] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_27b4_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l132_c21_9d89_return_output;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_e7fe] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_e7fe_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6486] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6486_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_61d2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_61d2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_8f00] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_8f00_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4669] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4669_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_8e6c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output;

     -- Submodule level 13
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_8e6c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6eed] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- Submodule level 14
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6eed_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_001b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- Submodule level 15
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_001b_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_302c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_d7f4] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- Submodule level 16
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_302c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_d7f4_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_c84f] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output;

     -- Submodule level 17
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c84f_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_b299] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- Submodule level 18
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_b299_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_683c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_8e84] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- Submodule level 19
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_8e84_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_683c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_3_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_c4ed] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_42ab] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- Submodule level 20
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_c4ed_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_42ab_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_4_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_6a38] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output;

     -- Submodule level 21
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_6a38_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_2_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_91bb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_54d5] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_fc1c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output;

     -- Submodule level 22
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_fc1c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_54d5_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_91bb_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_3_low_poly1305_h_l133_c13_3a49;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l132_c21_9d89] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_4553] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_353b] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- Submodule level 23
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_4553_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_353b_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l132_c21_9d89_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_1_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX[poly1305_h_l134_c22_74a0] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_cond;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iftrue;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_a9da] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output;

     -- Submodule level 24
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_a9da_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_MUX_poly1305_h_l134_c22_74a0_return_output;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_2_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_d037] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output;

     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- Submodule level 25
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_d037_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_high_poly1305_h_l134_c13_c226;
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_6e6c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output;

     -- Submodule level 26
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_6e6c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_1_low_poly1305_h_l133_c13_3a49;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_78a7] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output;

     -- Submodule level 27
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_78a7_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left := VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l131_c13_59af;
     -- FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_38af] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_left;
     FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right <= VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output := FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output;

     -- Submodule level 28
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49 := resize(VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_38af_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_3224] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_3224_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_0_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49,
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_1_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49,
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_2_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49,
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_3_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49,
     VAR_FOR_poly1305_h_l120_c5_7df6_ITER_4_FOR_poly1305_h_l123_c9_dbcd_ITER_0_low_poly1305_h_l133_c13_3a49);

     -- Submodule level 29
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_3224_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
