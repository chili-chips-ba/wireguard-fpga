-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 27
entity chacha20_block_0CLK_f1a496f6 is
port(
 state : in chacha20_state;
 return_output : out chacha20_state);
end chacha20_block_0CLK_f1a496f6;
architecture arch of chacha20_block_0CLK_f1a496f6 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- chacha20_block_step[chacha20_h_l72_c28_e45e]
signal chacha20_block_step_chacha20_h_l72_c28_e45e_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l72_c28_e45e_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l73_c28_04d0]
signal chacha20_block_step_chacha20_h_l73_c28_04d0_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l73_c28_04d0_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l74_c28_811c]
signal chacha20_block_step_chacha20_h_l74_c28_811c_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l74_c28_811c_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l75_c28_d3ec]
signal chacha20_block_step_chacha20_h_l75_c28_d3ec_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l76_c28_b3fd]
signal chacha20_block_step_chacha20_h_l76_c28_b3fd_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l77_c28_3088]
signal chacha20_block_step_chacha20_h_l77_c28_3088_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l77_c28_3088_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l78_c28_a4e0]
signal chacha20_block_step_chacha20_h_l78_c28_a4e0_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l79_c28_3e76]
signal chacha20_block_step_chacha20_h_l79_c28_3e76_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l79_c28_3e76_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l80_c28_e5e1]
signal chacha20_block_step_chacha20_h_l80_c28_e5e1_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output : chacha20_state;

-- chacha20_block_step[chacha20_h_l81_c29_93d8]
signal chacha20_block_step_chacha20_h_l81_c29_93d8_state0 : chacha20_state;
signal chacha20_block_step_chacha20_h_l81_c29_93d8_return_output : chacha20_state;

-- FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_a26c]
signal FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
signal FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);

function CONST_REF_RD_chacha20_state_chacha20_state_23da( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return chacha20_state is
 
  variable base : chacha20_state; 
  variable return_output : chacha20_state;
begin
      base.state(0) := ref_toks_0;
      base.state(1) := ref_toks_1;
      base.state(2) := ref_toks_2;
      base.state(3) := ref_toks_3;
      base.state(4) := ref_toks_4;
      base.state(5) := ref_toks_5;
      base.state(6) := ref_toks_6;
      base.state(7) := ref_toks_7;
      base.state(8) := ref_toks_8;
      base.state(9) := ref_toks_9;
      base.state(10) := ref_toks_10;
      base.state(11) := ref_toks_11;
      base.state(12) := ref_toks_12;
      base.state(13) := ref_toks_13;
      base.state(14) := ref_toks_14;
      base.state(15) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- chacha20_block_step_chacha20_h_l72_c28_e45e : 0 clocks latency
chacha20_block_step_chacha20_h_l72_c28_e45e : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l72_c28_e45e_state0,
chacha20_block_step_chacha20_h_l72_c28_e45e_return_output);

-- chacha20_block_step_chacha20_h_l73_c28_04d0 : 0 clocks latency
chacha20_block_step_chacha20_h_l73_c28_04d0 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l73_c28_04d0_state0,
chacha20_block_step_chacha20_h_l73_c28_04d0_return_output);

-- chacha20_block_step_chacha20_h_l74_c28_811c : 0 clocks latency
chacha20_block_step_chacha20_h_l74_c28_811c : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l74_c28_811c_state0,
chacha20_block_step_chacha20_h_l74_c28_811c_return_output);

-- chacha20_block_step_chacha20_h_l75_c28_d3ec : 0 clocks latency
chacha20_block_step_chacha20_h_l75_c28_d3ec : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l75_c28_d3ec_state0,
chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output);

-- chacha20_block_step_chacha20_h_l76_c28_b3fd : 0 clocks latency
chacha20_block_step_chacha20_h_l76_c28_b3fd : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l76_c28_b3fd_state0,
chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output);

-- chacha20_block_step_chacha20_h_l77_c28_3088 : 0 clocks latency
chacha20_block_step_chacha20_h_l77_c28_3088 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l77_c28_3088_state0,
chacha20_block_step_chacha20_h_l77_c28_3088_return_output);

-- chacha20_block_step_chacha20_h_l78_c28_a4e0 : 0 clocks latency
chacha20_block_step_chacha20_h_l78_c28_a4e0 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l78_c28_a4e0_state0,
chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output);

-- chacha20_block_step_chacha20_h_l79_c28_3e76 : 0 clocks latency
chacha20_block_step_chacha20_h_l79_c28_3e76 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l79_c28_3e76_state0,
chacha20_block_step_chacha20_h_l79_c28_3e76_return_output);

-- chacha20_block_step_chacha20_h_l80_c28_e5e1 : 0 clocks latency
chacha20_block_step_chacha20_h_l80_c28_e5e1 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l80_c28_e5e1_state0,
chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output);

-- chacha20_block_step_chacha20_h_l81_c29_93d8 : 0 clocks latency
chacha20_block_step_chacha20_h_l81_c29_93d8 : entity work.chacha20_block_step_0CLK_1e73dead port map (
chacha20_block_step_chacha20_h_l81_c29_93d8_state0,
chacha20_block_step_chacha20_h_l81_c29_93d8_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);

-- FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : 0 clocks latency
FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c : entity work.BIN_OP_PLUS_uint32_t_uint32_t_0CLK_de264c78 port map (
FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left,
FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right,
FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 state,
 -- All submodule outputs
 chacha20_block_step_chacha20_h_l72_c28_e45e_return_output,
 chacha20_block_step_chacha20_h_l73_c28_04d0_return_output,
 chacha20_block_step_chacha20_h_l74_c28_811c_return_output,
 chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output,
 chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output,
 chacha20_block_step_chacha20_h_l77_c28_3088_return_output,
 chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output,
 chacha20_block_step_chacha20_h_l79_c28_3e76_return_output,
 chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output,
 chacha20_block_step_chacha20_h_l81_c29_93d8_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output,
 FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : chacha20_state;
 variable VAR_state : chacha20_state;
 variable VAR_output : chacha20_state;
 variable VAR_step1 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_return_output : chacha20_state;
 variable VAR_step2 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_return_output : chacha20_state;
 variable VAR_step3 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_811c_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l74_c28_811c_return_output : chacha20_state;
 variable VAR_step4 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output : chacha20_state;
 variable VAR_step5 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output : chacha20_state;
 variable VAR_step6 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_3088_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l77_c28_3088_return_output : chacha20_state;
 variable VAR_step7 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output : chacha20_state;
 variable VAR_step8 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_return_output : chacha20_state;
 variable VAR_step9 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output : chacha20_state;
 variable VAR_step10 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_state0 : chacha20_state;
 variable VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output : chacha20_state;
 variable VAR_i : unsigned(3 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_output_state_0_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_output_state_1_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_output_state_2_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_output_state_3_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_output_state_4_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_output_state_5_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_output_state_6_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_output_state_7_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_output_state_8_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_output_state_9_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_output_state_10_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_output_state_11_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_output_state_12_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_output_state_13_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_output_state_14_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_output_state_15_chacha20_h_l87_c9_cff9 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_cc40_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_48bb_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_a4b6_return_output : chacha20_state;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_state := state;

     -- Submodule level 0
     VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_state0 := VAR_state;
     -- FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(5);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(0);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(15);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(3);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(13);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(7);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(11);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(9);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(8);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(4);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(2);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(12);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(6);

     -- chacha20_block_step[chacha20_h_l72_c28_e45e] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l72_c28_e45e_state0 <= VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_return_output := chacha20_block_step_chacha20_h_l72_c28_e45e_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(14);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(10);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c45_48bb] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_48bb_return_output := VAR_state.state(1);

     -- Submodule level 1
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c45_48bb_return_output;
     VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_state0 := VAR_chacha20_block_step_chacha20_h_l72_c28_e45e_return_output;
     -- chacha20_block_step[chacha20_h_l73_c28_04d0] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l73_c28_04d0_state0 <= VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_return_output := chacha20_block_step_chacha20_h_l73_c28_04d0_return_output;

     -- Submodule level 2
     VAR_chacha20_block_step_chacha20_h_l74_c28_811c_state0 := VAR_chacha20_block_step_chacha20_h_l73_c28_04d0_return_output;
     -- chacha20_block_step[chacha20_h_l74_c28_811c] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l74_c28_811c_state0 <= VAR_chacha20_block_step_chacha20_h_l74_c28_811c_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l74_c28_811c_return_output := chacha20_block_step_chacha20_h_l74_c28_811c_return_output;

     -- Submodule level 3
     VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_state0 := VAR_chacha20_block_step_chacha20_h_l74_c28_811c_return_output;
     -- chacha20_block_step[chacha20_h_l75_c28_d3ec] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l75_c28_d3ec_state0 <= VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output := chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output;

     -- Submodule level 4
     VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_state0 := VAR_chacha20_block_step_chacha20_h_l75_c28_d3ec_return_output;
     -- chacha20_block_step[chacha20_h_l76_c28_b3fd] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l76_c28_b3fd_state0 <= VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output := chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output;

     -- Submodule level 5
     VAR_chacha20_block_step_chacha20_h_l77_c28_3088_state0 := VAR_chacha20_block_step_chacha20_h_l76_c28_b3fd_return_output;
     -- chacha20_block_step[chacha20_h_l77_c28_3088] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l77_c28_3088_state0 <= VAR_chacha20_block_step_chacha20_h_l77_c28_3088_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l77_c28_3088_return_output := chacha20_block_step_chacha20_h_l77_c28_3088_return_output;

     -- Submodule level 6
     VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_state0 := VAR_chacha20_block_step_chacha20_h_l77_c28_3088_return_output;
     -- chacha20_block_step[chacha20_h_l78_c28_a4e0] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l78_c28_a4e0_state0 <= VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output := chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output;

     -- Submodule level 7
     VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_state0 := VAR_chacha20_block_step_chacha20_h_l78_c28_a4e0_return_output;
     -- chacha20_block_step[chacha20_h_l79_c28_3e76] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l79_c28_3e76_state0 <= VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_return_output := chacha20_block_step_chacha20_h_l79_c28_3e76_return_output;

     -- Submodule level 8
     VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_state0 := VAR_chacha20_block_step_chacha20_h_l79_c28_3e76_return_output;
     -- chacha20_block_step[chacha20_h_l80_c28_e5e1] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l80_c28_e5e1_state0 <= VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output := chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output;

     -- Submodule level 9
     VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_state0 := VAR_chacha20_block_step_chacha20_h_l80_c28_e5e1_return_output;
     -- chacha20_block_step[chacha20_h_l81_c29_93d8] LATENCY=0
     -- Inputs
     chacha20_block_step_chacha20_h_l81_c29_93d8_state0 <= VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_state0;
     -- Outputs
     VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output := chacha20_block_step_chacha20_h_l81_c29_93d8_return_output;

     -- Submodule level 10
     -- FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(5);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(9);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(11);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(15);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(0);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(3);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(10);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(6);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(12);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(14);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(2);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(4);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(1);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(13);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(7);

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_h_l87_c27_cc40] LATENCY=0
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_cc40_return_output := VAR_chacha20_block_step_chacha20_h_l81_c29_93d8_return_output.state(8);

     -- Submodule level 11
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_h_l87_c27_cc40_return_output;
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left := VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_h_l87_c27_cc40_return_output;
     -- FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS[chacha20_h_l87_c27_a26c] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_left;
     FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right <= VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_right;
     -- Outputs
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output := FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output;

     -- Submodule level 12
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_output_state_0_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_output_state_10_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_output_state_11_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_output_state_12_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_output_state_13_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_output_state_14_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_output_state_15_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_output_state_1_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_output_state_2_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_output_state_3_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_output_state_4_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_output_state_5_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_output_state_6_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_output_state_7_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_output_state_8_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_output_state_9_chacha20_h_l87_c9_cff9 := resize(VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_BIN_OP_PLUS_chacha20_h_l87_c27_a26c_return_output, 32);
     -- CONST_REF_RD_chacha20_state_chacha20_state_23da[chacha20_h_l90_c12_a4b6] LATENCY=0
     VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_a4b6_return_output := CONST_REF_RD_chacha20_state_chacha20_state_23da(
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_0_output_state_0_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_1_output_state_1_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_2_output_state_2_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_3_output_state_3_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_4_output_state_4_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_5_output_state_5_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_6_output_state_6_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_7_output_state_7_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_8_output_state_8_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_9_output_state_9_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_10_output_state_10_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_11_output_state_11_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_12_output_state_12_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_13_output_state_13_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_14_output_state_14_chacha20_h_l87_c9_cff9,
     VAR_FOR_chacha20_h_l85_c5_2cc3_ITER_15_output_state_15_chacha20_h_l87_c9_cff9);

     -- Submodule level 13
     VAR_return_output := VAR_CONST_REF_RD_chacha20_state_chacha20_state_23da_chacha20_h_l90_c12_a4b6_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
