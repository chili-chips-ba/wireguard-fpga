-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.01818181818181818, 0.03636363636363636, 0.054545454545454536, 0.07272727272727272, 0.09090909090909093, 0.1090909090909091, 0.1272727272727273, 0.14545454545454548, 0.16363636363636366, 0.18181818181818185, 0.20000000000000004, 0.21818181818181823, 0.23636363636363641, 0.2545454545454546, 0.27272727272727276, 0.29090909090909095, 0.30909090909090914, 0.3272727272727273, 0.3454545454545455, 0.3636363636363637, 0.38181818181818195, 0.4000000000000001, 0.41818181818181827, 0.43636363636363645, 0.45454545454545464, 0.47272727272727283, 0.49090909090909096, 0.5090909090909091, 0.5272727272727273, 0.5454545454545455, 0.5636363636363637, 0.5818181818181819, 0.6000000000000001, 0.6181818181818183, 0.6363636363636365, 0.6545454545454547, 0.6727272727272728, 0.690909090909091, 0.7090909090909092, 0.7272727272727274, 0.7454545454545455, 0.7636363636363639, 0.7818181818181821, 0.8000000000000002, 0.8181818181818183, 0.8363636363636365, 0.8545454545454547, 0.8727272727272729, 0.8909090909090911, 0.9090909090909093, 0.9272727272727275, 0.9454545454545457, 0.9636363636363638, 0.9818181818181819]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 69
entity chacha20_decrypt_loop_body_54CLK_0d2f63f1 is
port(
 clk : in std_logic;
 inputs : in chacha20_decrypt_loop_body_in_t;
 return_output : out axis512_t);
end chacha20_decrypt_loop_body_54CLK_0d2f63f1;
architecture arch of chacha20_decrypt_loop_body_54CLK_0d2f63f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 54;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 1
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 2
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 3
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 4
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 5
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 6
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 7
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 8
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 9
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 10
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 11
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 12
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 13
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 14
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 15
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 16
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 17
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 18
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 19
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 20
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 21
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 22
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 23
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 24
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 25
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 26
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 27
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 28
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 29
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 30
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 31
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 32
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 33
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 34
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 35
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 36
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 37
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 38
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 39
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 40
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 41
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 42
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 43
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 44
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 45
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 46
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 47
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 48
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 49
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 50
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 51
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 52
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Stage 53
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal REG_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal COMB_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
-- Each function instance gets signals
-- chacha20_init[chacha20_h_l216_c26_71b5]
signal chacha20_init_chacha20_h_l216_c26_71b5_key : uint8_t_32;
signal chacha20_init_chacha20_h_l216_c26_71b5_nonce : uint8_t_12;
signal chacha20_init_chacha20_h_l216_c26_71b5_counter : unsigned(31 downto 0);
signal chacha20_init_chacha20_h_l216_c26_71b5_return_output : chacha20_state;

-- chacha20_block[chacha20_h_l217_c26_8f03]
signal chacha20_block_chacha20_h_l217_c26_8f03_state : chacha20_state;
signal chacha20_block_chacha20_h_l217_c26_8f03_return_output : chacha20_state;

-- chacha20_state_to_bytes[chacha20_h_l220_c38_26de]
signal chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x : chacha20_state;
signal chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output : uint8_t_array_64_t;

-- FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

-- FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR[chacha20_h_l228_c19_168d]
signal FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
signal FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_64_uint8_t_64_62ba( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned) return uint8_t_64 is
 
  variable base : uint8_t_64; 
  variable return_output : uint8_t_64;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;
      base(12) := ref_toks_12;
      base(13) := ref_toks_13;
      base(14) := ref_toks_14;
      base(15) := ref_toks_15;
      base(16) := ref_toks_16;
      base(17) := ref_toks_17;
      base(18) := ref_toks_18;
      base(19) := ref_toks_19;
      base(20) := ref_toks_20;
      base(21) := ref_toks_21;
      base(22) := ref_toks_22;
      base(23) := ref_toks_23;
      base(24) := ref_toks_24;
      base(25) := ref_toks_25;
      base(26) := ref_toks_26;
      base(27) := ref_toks_27;
      base(28) := ref_toks_28;
      base(29) := ref_toks_29;
      base(30) := ref_toks_30;
      base(31) := ref_toks_31;
      base(32) := ref_toks_32;
      base(33) := ref_toks_33;
      base(34) := ref_toks_34;
      base(35) := ref_toks_35;
      base(36) := ref_toks_36;
      base(37) := ref_toks_37;
      base(38) := ref_toks_38;
      base(39) := ref_toks_39;
      base(40) := ref_toks_40;
      base(41) := ref_toks_41;
      base(42) := ref_toks_42;
      base(43) := ref_toks_43;
      base(44) := ref_toks_44;
      base(45) := ref_toks_45;
      base(46) := ref_toks_46;
      base(47) := ref_toks_47;
      base(48) := ref_toks_48;
      base(49) := ref_toks_49;
      base(50) := ref_toks_50;
      base(51) := ref_toks_51;
      base(52) := ref_toks_52;
      base(53) := ref_toks_53;
      base(54) := ref_toks_54;
      base(55) := ref_toks_55;
      base(56) := ref_toks_56;
      base(57) := ref_toks_57;
      base(58) := ref_toks_58;
      base(59) := ref_toks_59;
      base(60) := ref_toks_60;
      base(61) := ref_toks_61;
      base(62) := ref_toks_62;
      base(63) := ref_toks_63;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis512_t_axis512_t_774e( ref_toks_0 : axis512_t;
 ref_toks_1 : uint8_t_64) return axis512_t is
 
  variable base : axis512_t; 
  variable return_output : axis512_t;
begin
      base := ref_toks_0;
      base.tdata := ref_toks_1;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- chacha20_init_chacha20_h_l216_c26_71b5 : 0 clocks latency
chacha20_init_chacha20_h_l216_c26_71b5 : entity work.chacha20_init_0CLK_50a1b8d0 port map (
chacha20_init_chacha20_h_l216_c26_71b5_key,
chacha20_init_chacha20_h_l216_c26_71b5_nonce,
chacha20_init_chacha20_h_l216_c26_71b5_counter,
chacha20_init_chacha20_h_l216_c26_71b5_return_output);

-- chacha20_block_chacha20_h_l217_c26_8f03 : 54 clocks latency
chacha20_block_chacha20_h_l217_c26_8f03 : entity work.chacha20_block_54CLK_608c4823 port map (
clk,
chacha20_block_chacha20_h_l217_c26_8f03_state,
chacha20_block_chacha20_h_l217_c26_8f03_return_output);

-- chacha20_state_to_bytes_chacha20_h_l220_c38_26de : 0 clocks latency
chacha20_state_to_bytes_chacha20_h_l220_c38_26de : entity work.chacha20_state_to_bytes_0CLK_d3fba2d7 port map (
chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x,
chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

-- FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d : 0 clocks latency
FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right,
FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 inputs,
 -- Registers
 -- Stage 0
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 1
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 2
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 3
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 4
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 5
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 6
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 7
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 8
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 9
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 10
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 11
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 12
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 13
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 14
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 15
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 16
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 17
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 18
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 19
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 20
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 21
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 22
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 23
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 24
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 25
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 26
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 27
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 28
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 29
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 30
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 31
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 32
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 33
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 34
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 35
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 36
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 37
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 38
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 39
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 40
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 41
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 42
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 43
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 44
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 45
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 46
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 47
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 48
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 49
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 50
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 51
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 52
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- Stage 53
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left,
 REG_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
 -- All submodule outputs
 chacha20_init_chacha20_h_l216_c26_71b5_return_output,
 chacha20_block_chacha20_h_l217_c26_8f03_return_output,
 chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
 FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis512_t;
 variable VAR_inputs : chacha20_decrypt_loop_body_in_t;
 variable VAR_in_data : uint8_t_64;
 variable VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output : uint8_t_64;
 variable VAR_key : uint8_t_32;
 variable VAR_CONST_REF_RD_uint8_t_32_chacha20_decrypt_loop_body_in_t_key_d41d_chacha20_h_l212_c21_05d4_return_output : uint8_t_32;
 variable VAR_nonce : uint8_t_12;
 variable VAR_CONST_REF_RD_uint8_t_12_chacha20_decrypt_loop_body_in_t_nonce_d41d_chacha20_h_l213_c23_dcf4_return_output : uint8_t_12;
 variable VAR_counter : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint32_t_chacha20_decrypt_loop_body_in_t_counter_d41d_chacha20_h_l214_c22_73ac_return_output : unsigned(31 downto 0);
 variable VAR_state : chacha20_state;
 variable VAR_chacha20_init_chacha20_h_l216_c26_71b5_key : uint8_t_32;
 variable VAR_chacha20_init_chacha20_h_l216_c26_71b5_nonce : uint8_t_12;
 variable VAR_chacha20_init_chacha20_h_l216_c26_71b5_counter : unsigned(31 downto 0);
 variable VAR_chacha20_init_chacha20_h_l216_c26_71b5_return_output : chacha20_state;
 variable VAR_block : chacha20_state;
 variable VAR_chacha20_block_chacha20_h_l217_c26_8f03_state : chacha20_state;
 variable VAR_chacha20_block_chacha20_h_l217_c26_8f03_return_output : chacha20_state;
 variable VAR_block_bytes_t : uint8_t_array_64_t;
 variable VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x : chacha20_state;
 variable VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output : uint8_t_array_64_t;
 variable VAR_block_bytes : uint8_t_64;
 variable VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output : uint8_t_64;
 variable VAR_out_data : uint8_t_64;
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c19_594b_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c32_44b5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output : unsigned(7 downto 0);
 variable VAR_axis_out : axis512_t;
 variable VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output : axis512_t;
 variable VAR_CONST_REF_RD_uint8_t_64_uint8_t_64_62ba_chacha20_h_l233_c20_5d4d_return_output : uint8_t_64;
 variable VAR_CONST_REF_RD_axis512_t_axis512_t_774e_chacha20_h_l234_c10_0437_return_output : axis512_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_inputs := inputs;

     -- Submodule level 0
     -- CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d[chacha20_h_l231_c24_0fd7] LATENCY=0
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := VAR_inputs.axis_in;

     -- CONST_REF_RD_uint32_t_chacha20_decrypt_loop_body_in_t_counter_d41d[chacha20_h_l214_c22_73ac] LATENCY=0
     VAR_CONST_REF_RD_uint32_t_chacha20_decrypt_loop_body_in_t_counter_d41d_chacha20_h_l214_c22_73ac_return_output := VAR_inputs.counter;

     -- CONST_REF_RD_uint8_t_12_chacha20_decrypt_loop_body_in_t_nonce_d41d[chacha20_h_l213_c23_dcf4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_12_chacha20_decrypt_loop_body_in_t_nonce_d41d_chacha20_h_l213_c23_dcf4_return_output := VAR_inputs.nonce;

     -- CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d[chacha20_h_l211_c25_87c0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output := VAR_inputs.axis_in.tdata;

     -- CONST_REF_RD_uint8_t_32_chacha20_decrypt_loop_body_in_t_key_d41d[chacha20_h_l212_c21_05d4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_32_chacha20_decrypt_loop_body_in_t_key_d41d_chacha20_h_l212_c21_05d4_return_output := VAR_inputs.key;

     -- Submodule level 1
     VAR_chacha20_init_chacha20_h_l216_c26_71b5_counter := VAR_CONST_REF_RD_uint32_t_chacha20_decrypt_loop_body_in_t_counter_d41d_chacha20_h_l214_c22_73ac_return_output;
     VAR_chacha20_init_chacha20_h_l216_c26_71b5_nonce := VAR_CONST_REF_RD_uint8_t_12_chacha20_decrypt_loop_body_in_t_nonce_d41d_chacha20_h_l213_c23_dcf4_return_output;
     VAR_chacha20_init_chacha20_h_l216_c26_71b5_key := VAR_CONST_REF_RD_uint8_t_32_chacha20_decrypt_loop_body_in_t_key_d41d_chacha20_h_l212_c21_05d4_return_output;
     -- FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(48);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(20);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(27);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(59);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(45);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(46);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(41);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(53);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(6);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(47);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(56);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(63);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(10);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(61);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(2);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(43);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(23);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(40);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(25);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(49);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(9);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(4);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(5);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(52);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(60);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(12);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(3);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(30);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(21);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(32);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(29);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(44);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(58);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(55);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(34);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(36);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(24);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(0);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(57);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(1);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(11);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(18);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(17);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(14);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(13);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(7);

     -- chacha20_init[chacha20_h_l216_c26_71b5] LATENCY=0
     -- Inputs
     chacha20_init_chacha20_h_l216_c26_71b5_key <= VAR_chacha20_init_chacha20_h_l216_c26_71b5_key;
     chacha20_init_chacha20_h_l216_c26_71b5_nonce <= VAR_chacha20_init_chacha20_h_l216_c26_71b5_nonce;
     chacha20_init_chacha20_h_l216_c26_71b5_counter <= VAR_chacha20_init_chacha20_h_l216_c26_71b5_counter;
     -- Outputs
     VAR_chacha20_init_chacha20_h_l216_c26_71b5_return_output := chacha20_init_chacha20_h_l216_c26_71b5_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(35);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(28);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(19);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(38);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(50);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(33);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(54);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(8);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(62);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(39);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(51);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(22);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(15);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(31);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(42);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(37);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(26);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d[chacha20_h_l228_c19_594b] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c19_594b_return_output := VAR_CONST_REF_RD_uint8_t_64_chacha20_decrypt_loop_body_in_t_axis_in_tdata_d41d_chacha20_h_l211_c25_87c0_return_output(16);

     -- Submodule level 2
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c19_594b_return_output;
     VAR_chacha20_block_chacha20_h_l217_c26_8f03_state := VAR_chacha20_init_chacha20_h_l216_c26_71b5_return_output;
     -- chacha20_block[chacha20_h_l217_c26_8f03] LATENCY=54
     -- Inputs
     chacha20_block_chacha20_h_l217_c26_8f03_state <= VAR_chacha20_block_chacha20_h_l217_c26_8f03_state;

     -- Write to comb signals
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 26 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 27 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 28 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 29 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 30 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 31 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 32 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 33 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 34 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 35 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 36 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 37 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 38 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 39 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 40 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 41 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 42 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 43 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 44 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 45 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 46 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 47 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 48 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 49 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 50 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 51 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 52 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 53 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;

     -- Write to comb signals
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     COMB_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
   elsif STAGE = 54 then
     -- Read from prev stage
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left := REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output := REG_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Submodule outputs
     VAR_chacha20_block_chacha20_h_l217_c26_8f03_return_output := chacha20_block_chacha20_h_l217_c26_8f03_return_output;

     -- Submodule level 0
     VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x := VAR_chacha20_block_chacha20_h_l217_c26_8f03_return_output;
     -- chacha20_state_to_bytes[chacha20_h_l220_c38_26de] LATENCY=0
     -- Inputs
     chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x <= VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_x;
     -- Outputs
     VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output := chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d[chacha20_h_l221_c29_09c2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output := VAR_chacha20_state_to_bytes_chacha20_h_l220_c38_26de_return_output.data;

     -- Submodule level 2
     -- FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(38);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(52);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(30);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(54);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(26);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(33);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(24);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(40);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(15);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(62);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(42);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(41);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(61);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(22);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(29);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(27);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(35);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(46);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(23);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(39);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(58);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(34);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(1);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(28);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(3);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(7);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(11);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(37);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(59);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(47);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(49);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(16);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(10);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(51);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(60);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(9);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(14);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(55);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(17);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(45);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(36);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(31);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(5);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(44);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(12);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(53);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(32);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(8);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(20);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(2);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(56);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(0);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(18);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(21);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(4);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(6);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(43);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(63);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(13);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(57);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(19);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(50);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(48);

     -- FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d[chacha20_h_l228_c32_44b5] LATENCY=0
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c32_44b5_return_output := VAR_CONST_REF_RD_uint8_t_64_uint8_t_array_64_t_data_d41d_chacha20_h_l221_c29_09c2_return_output(25);

     -- Submodule level 3
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_CONST_REF_RD_uint8_t_uint8_t_64_0_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_CONST_REF_RD_uint8_t_uint8_t_64_10_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_CONST_REF_RD_uint8_t_uint8_t_64_11_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_CONST_REF_RD_uint8_t_uint8_t_64_12_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_CONST_REF_RD_uint8_t_uint8_t_64_13_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_CONST_REF_RD_uint8_t_uint8_t_64_14_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_CONST_REF_RD_uint8_t_uint8_t_64_15_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_CONST_REF_RD_uint8_t_uint8_t_64_16_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_CONST_REF_RD_uint8_t_uint8_t_64_17_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_CONST_REF_RD_uint8_t_uint8_t_64_18_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_CONST_REF_RD_uint8_t_uint8_t_64_19_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_CONST_REF_RD_uint8_t_uint8_t_64_1_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_CONST_REF_RD_uint8_t_uint8_t_64_20_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_CONST_REF_RD_uint8_t_uint8_t_64_21_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_CONST_REF_RD_uint8_t_uint8_t_64_22_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_CONST_REF_RD_uint8_t_uint8_t_64_23_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_CONST_REF_RD_uint8_t_uint8_t_64_24_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_CONST_REF_RD_uint8_t_uint8_t_64_25_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_CONST_REF_RD_uint8_t_uint8_t_64_26_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_CONST_REF_RD_uint8_t_uint8_t_64_27_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_CONST_REF_RD_uint8_t_uint8_t_64_28_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_CONST_REF_RD_uint8_t_uint8_t_64_29_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_CONST_REF_RD_uint8_t_uint8_t_64_2_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_CONST_REF_RD_uint8_t_uint8_t_64_30_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_CONST_REF_RD_uint8_t_uint8_t_64_31_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_CONST_REF_RD_uint8_t_uint8_t_64_32_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_CONST_REF_RD_uint8_t_uint8_t_64_33_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_CONST_REF_RD_uint8_t_uint8_t_64_34_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_CONST_REF_RD_uint8_t_uint8_t_64_35_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_CONST_REF_RD_uint8_t_uint8_t_64_36_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_CONST_REF_RD_uint8_t_uint8_t_64_37_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_CONST_REF_RD_uint8_t_uint8_t_64_38_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_CONST_REF_RD_uint8_t_uint8_t_64_39_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_CONST_REF_RD_uint8_t_uint8_t_64_3_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_CONST_REF_RD_uint8_t_uint8_t_64_40_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_CONST_REF_RD_uint8_t_uint8_t_64_41_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_CONST_REF_RD_uint8_t_uint8_t_64_42_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_CONST_REF_RD_uint8_t_uint8_t_64_43_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_CONST_REF_RD_uint8_t_uint8_t_64_44_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_CONST_REF_RD_uint8_t_uint8_t_64_45_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_CONST_REF_RD_uint8_t_uint8_t_64_46_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_CONST_REF_RD_uint8_t_uint8_t_64_47_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_CONST_REF_RD_uint8_t_uint8_t_64_48_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_CONST_REF_RD_uint8_t_uint8_t_64_49_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_CONST_REF_RD_uint8_t_uint8_t_64_4_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_CONST_REF_RD_uint8_t_uint8_t_64_50_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_CONST_REF_RD_uint8_t_uint8_t_64_51_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_CONST_REF_RD_uint8_t_uint8_t_64_52_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_CONST_REF_RD_uint8_t_uint8_t_64_53_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_CONST_REF_RD_uint8_t_uint8_t_64_54_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_CONST_REF_RD_uint8_t_uint8_t_64_55_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_CONST_REF_RD_uint8_t_uint8_t_64_56_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_CONST_REF_RD_uint8_t_uint8_t_64_57_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_CONST_REF_RD_uint8_t_uint8_t_64_58_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_CONST_REF_RD_uint8_t_uint8_t_64_59_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_CONST_REF_RD_uint8_t_uint8_t_64_5_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_CONST_REF_RD_uint8_t_uint8_t_64_60_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_CONST_REF_RD_uint8_t_uint8_t_64_61_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_CONST_REF_RD_uint8_t_uint8_t_64_62_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_CONST_REF_RD_uint8_t_uint8_t_64_63_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_CONST_REF_RD_uint8_t_uint8_t_64_6_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_CONST_REF_RD_uint8_t_uint8_t_64_7_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_CONST_REF_RD_uint8_t_uint8_t_64_8_d41d_chacha20_h_l228_c32_44b5_return_output;
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right := VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_CONST_REF_RD_uint8_t_uint8_t_64_9_d41d_chacha20_h_l228_c32_44b5_return_output;
     -- FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR[chacha20_h_l228_c19_168d] LATENCY=0
     -- Inputs
     FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right <= VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_right;
     -- Outputs
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output := FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output;

     -- Submodule level 4
     -- CONST_REF_RD_uint8_t_64_uint8_t_64_62ba[chacha20_h_l233_c20_5d4d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_64_uint8_t_64_62ba_chacha20_h_l233_c20_5d4d_return_output := CONST_REF_RD_uint8_t_64_uint8_t_64_62ba(
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output,
     VAR_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_return_output);

     -- Submodule level 5
     -- CONST_REF_RD_axis512_t_axis512_t_774e[chacha20_h_l234_c10_0437] LATENCY=0
     VAR_CONST_REF_RD_axis512_t_axis512_t_774e_chacha20_h_l234_c10_0437_return_output := CONST_REF_RD_axis512_t_axis512_t_774e(
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output,
     VAR_CONST_REF_RD_uint8_t_64_uint8_t_64_62ba_chacha20_h_l233_c20_5d4d_return_output);

     -- Submodule level 6
     VAR_return_output := VAR_CONST_REF_RD_axis512_t_axis512_t_774e_chacha20_h_l234_c10_0437_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE0_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE0_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 1
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE1_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE1_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 2
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE2_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE2_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 3
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE3_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE3_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 4
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE4_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE4_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 5
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE5_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE5_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 6
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE6_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE6_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 7
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE7_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE7_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 8
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE8_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE8_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 9
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE9_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE9_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 10
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE10_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE10_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 11
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE11_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE11_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 12
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE12_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE12_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 13
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE13_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE13_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 14
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE14_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE14_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 15
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE15_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE15_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 16
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE16_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE16_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 17
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE17_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE17_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 18
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE18_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE18_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 19
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE19_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE19_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 20
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE20_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE20_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 21
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE21_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE21_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 22
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE22_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE22_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 23
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE23_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE23_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 24
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE24_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE24_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 25
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE25_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE25_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 26
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE26_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE26_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 27
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE27_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE27_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 28
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE28_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE28_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 29
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE29_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE29_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 30
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE30_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE30_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 31
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE31_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE31_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 32
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE32_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE32_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 33
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE33_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE33_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 34
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE34_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE34_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 35
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE35_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE35_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 36
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE36_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE36_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 37
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE37_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE37_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 38
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE38_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE38_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 39
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE39_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE39_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 40
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE40_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE40_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 41
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE41_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE41_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 42
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE42_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE42_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 43
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE43_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE43_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 44
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE44_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE44_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 45
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE45_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE45_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 46
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE46_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE46_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 47
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE47_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE47_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 48
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE48_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE48_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 49
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE49_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE49_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 50
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE50_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE50_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 51
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE51_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE51_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 52
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE52_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE52_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
     -- Stage 53
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_0_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_1_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_2_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_3_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_4_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_5_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_6_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_7_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_8_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_9_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_10_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_11_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_12_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_13_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_14_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_15_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_16_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_17_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_18_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_19_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_20_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_21_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_22_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_23_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_24_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_25_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_26_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_27_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_28_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_29_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_30_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_31_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_32_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_33_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_34_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_35_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_36_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_37_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_38_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_39_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_40_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_41_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_42_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_43_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_44_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_45_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_46_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_47_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_48_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_49_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_50_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_51_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_52_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_53_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_54_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_55_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_56_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_57_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_58_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_59_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_60_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_61_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_62_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left <= COMB_STAGE53_FOR_chacha20_h_l226_c3_2e21_ITER_63_BIN_OP_XOR_chacha20_h_l228_c19_168d_left;
     REG_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output <= COMB_STAGE53_CONST_REF_RD_axis512_t_chacha20_decrypt_loop_body_in_t_axis_in_d41d_chacha20_h_l231_c24_0fd7_return_output;
 end if;
end process;

end arch;
