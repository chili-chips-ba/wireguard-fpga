mem['h0000] = 32'h00001517;
mem['h0001] = 32'h18050513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h00418593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h0E0000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'hFE010113;
mem['h001D] = 32'h00A12623;
mem['h001E] = 32'h0001A783;
mem['h001F] = 32'h00078713;
mem['h0020] = 32'h100007B7;
mem['h0021] = 32'h00078793;
mem['h0022] = 32'h00F707B3;
mem['h0023] = 32'h00F12E23;
mem['h0024] = 32'h0001A703;
mem['h0025] = 32'h00C12783;
mem['h0026] = 32'h00F70733;
mem['h0027] = 32'h00E1A023;
mem['h0028] = 32'h0001A703;
mem['h0029] = 32'h000017B7;
mem['h002A] = 32'h80078793;
mem['h002B] = 32'h00E7D463;
mem['h002C] = 32'h00100073;
mem['h002D] = 32'h01C12783;
mem['h002E] = 32'h00078513;
mem['h002F] = 32'h02010113;
mem['h0030] = 32'h00008067;
mem['h0031] = 32'hFD010113;
mem['h0032] = 32'h02112623;
mem['h0033] = 32'h00A12623;
mem['h0034] = 32'h00C12783;
mem['h0035] = 32'h00078513;
mem['h0036] = 32'hF99FF0EF;
mem['h0037] = 32'h00A12E23;
mem['h0038] = 32'h01C12783;
mem['h0039] = 32'h00078513;
mem['h003A] = 32'h02C12083;
mem['h003B] = 32'h03010113;
mem['h003C] = 32'h00008067;
mem['h003D] = 32'hFF010113;
mem['h003E] = 32'h00A12623;
mem['h003F] = 32'h00000013;
mem['h0040] = 32'h01010113;
mem['h0041] = 32'h00008067;
mem['h0042] = 32'hFE010113;
mem['h0043] = 32'h00A12623;
mem['h0044] = 32'h00012E23;
mem['h0045] = 32'h0100006F;
mem['h0046] = 32'h01C12783;
mem['h0047] = 32'h00178793;
mem['h0048] = 32'h00F12E23;
mem['h0049] = 32'h01C12783;
mem['h004A] = 32'h00C12703;
mem['h004B] = 32'h00E7B7B3;
mem['h004C] = 32'h0FF7F793;
mem['h004D] = 32'hFE0792E3;
mem['h004E] = 32'h00000013;
mem['h004F] = 32'h00000013;
mem['h0050] = 32'h02010113;
mem['h0051] = 32'h00008067;
mem['h0052] = 32'hFC010113;
mem['h0053] = 32'h02112E23;
mem['h0054] = 32'h02812C23;
mem['h0055] = 32'h02400513;
mem['h0056] = 32'hF6DFF0EF;
mem['h0057] = 32'h00050793;
mem['h0058] = 32'h00078413;
mem['h0059] = 32'h200005B7;
mem['h005A] = 32'h00040513;
mem['h005B] = 32'h7D4000EF;
mem['h005C] = 32'h02812623;
mem['h005D] = 32'h000017B7;
mem['h005E] = 32'h06C78593;
mem['h005F] = 32'h02C12503;
mem['h0060] = 32'h205000EF;
mem['h0061] = 32'h02C12503;
mem['h0062] = 32'h351000EF;
mem['h0063] = 32'h00C10793;
mem['h0064] = 32'h00078593;
mem['h0065] = 32'h02C12503;
mem['h0066] = 32'h23D000EF;
mem['h0067] = 32'hFF1FF06F;
mem['h0068] = 32'hFF010113;
mem['h0069] = 32'h00A12623;
mem['h006A] = 32'h00B12423;
mem['h006B] = 32'h00C12783;
mem['h006C] = 32'h00812703;
mem['h006D] = 32'h00E7A023;
mem['h006E] = 32'h00000013;
mem['h006F] = 32'h01010113;
mem['h0070] = 32'h00008067;
mem['h0071] = 32'hFF010113;
mem['h0072] = 32'h00A12623;
mem['h0073] = 32'h00B12423;
mem['h0074] = 32'h00C12783;
mem['h0075] = 32'h00812703;
mem['h0076] = 32'h00E7A023;
mem['h0077] = 32'h00000013;
mem['h0078] = 32'h01010113;
mem['h0079] = 32'h00008067;
mem['h007A] = 32'hFF010113;
mem['h007B] = 32'h00A12623;
mem['h007C] = 32'h00B12423;
mem['h007D] = 32'h00C12783;
mem['h007E] = 32'h00812703;
mem['h007F] = 32'h00E7A023;
mem['h0080] = 32'h00000013;
mem['h0081] = 32'h01010113;
mem['h0082] = 32'h00008067;
mem['h0083] = 32'hFF010113;
mem['h0084] = 32'h00A12623;
mem['h0085] = 32'h00B12423;
mem['h0086] = 32'h00C12783;
mem['h0087] = 32'h00812703;
mem['h0088] = 32'h00E7A023;
mem['h0089] = 32'h00000013;
mem['h008A] = 32'h01010113;
mem['h008B] = 32'h00008067;
mem['h008C] = 32'hFF010113;
mem['h008D] = 32'h00A12623;
mem['h008E] = 32'h00B12423;
mem['h008F] = 32'h00C12783;
mem['h0090] = 32'h00812703;
mem['h0091] = 32'h00E7A023;
mem['h0092] = 32'h00000013;
mem['h0093] = 32'h01010113;
mem['h0094] = 32'h00008067;
mem['h0095] = 32'hFF010113;
mem['h0096] = 32'h00A12623;
mem['h0097] = 32'h00B12423;
mem['h0098] = 32'h00C12783;
mem['h0099] = 32'h00812703;
mem['h009A] = 32'h00E7A023;
mem['h009B] = 32'h00000013;
mem['h009C] = 32'h01010113;
mem['h009D] = 32'h00008067;
mem['h009E] = 32'hFF010113;
mem['h009F] = 32'h00A12623;
mem['h00A0] = 32'h00B12423;
mem['h00A1] = 32'h00C12783;
mem['h00A2] = 32'h00812703;
mem['h00A3] = 32'h00E7A023;
mem['h00A4] = 32'h00000013;
mem['h00A5] = 32'h01010113;
mem['h00A6] = 32'h00008067;
mem['h00A7] = 32'hFE010113;
mem['h00A8] = 32'h00112E23;
mem['h00A9] = 32'h00812C23;
mem['h00AA] = 32'h00A12623;
mem['h00AB] = 32'h00B12423;
mem['h00AC] = 32'h00400513;
mem['h00AD] = 32'hE11FF0EF;
mem['h00AE] = 32'h00050793;
mem['h00AF] = 32'h00078413;
mem['h00B0] = 32'h00812583;
mem['h00B1] = 32'h00040513;
mem['h00B2] = 32'hED9FF0EF;
mem['h00B3] = 32'h00C12783;
mem['h00B4] = 32'h0087A023;
mem['h00B5] = 32'h00400513;
mem['h00B6] = 32'hDEDFF0EF;
mem['h00B7] = 32'h00050793;
mem['h00B8] = 32'h00078413;
mem['h00B9] = 32'h00812783;
mem['h00BA] = 32'h00478793;
mem['h00BB] = 32'h00078593;
mem['h00BC] = 32'h00040513;
mem['h00BD] = 32'hED1FF0EF;
mem['h00BE] = 32'h00C12783;
mem['h00BF] = 32'h0087A223;
mem['h00C0] = 32'h00400513;
mem['h00C1] = 32'hDC1FF0EF;
mem['h00C2] = 32'h00050793;
mem['h00C3] = 32'h00078413;
mem['h00C4] = 32'h00812783;
mem['h00C5] = 32'h00878793;
mem['h00C6] = 32'h00078593;
mem['h00C7] = 32'h00040513;
mem['h00C8] = 32'hEC9FF0EF;
mem['h00C9] = 32'h00C12783;
mem['h00CA] = 32'h0087A423;
mem['h00CB] = 32'h00400513;
mem['h00CC] = 32'hD95FF0EF;
mem['h00CD] = 32'h00050793;
mem['h00CE] = 32'h00078413;
mem['h00CF] = 32'h00812783;
mem['h00D0] = 32'h00C78793;
mem['h00D1] = 32'h00078593;
mem['h00D2] = 32'h00040513;
mem['h00D3] = 32'hEC1FF0EF;
mem['h00D4] = 32'h00C12783;
mem['h00D5] = 32'h0087A623;
mem['h00D6] = 32'h00400513;
mem['h00D7] = 32'hD69FF0EF;
mem['h00D8] = 32'h00050793;
mem['h00D9] = 32'h00078413;
mem['h00DA] = 32'h00812783;
mem['h00DB] = 32'h01078793;
mem['h00DC] = 32'h00078593;
mem['h00DD] = 32'h00040513;
mem['h00DE] = 32'hEB9FF0EF;
mem['h00DF] = 32'h00C12783;
mem['h00E0] = 32'h0087A823;
mem['h00E1] = 32'h00400513;
mem['h00E2] = 32'hD3DFF0EF;
mem['h00E3] = 32'h00050793;
mem['h00E4] = 32'h00078413;
mem['h00E5] = 32'h00812783;
mem['h00E6] = 32'h01478793;
mem['h00E7] = 32'h00078593;
mem['h00E8] = 32'h00040513;
mem['h00E9] = 32'hEB1FF0EF;
mem['h00EA] = 32'h00C12783;
mem['h00EB] = 32'h0087AA23;
mem['h00EC] = 32'h00400513;
mem['h00ED] = 32'hD11FF0EF;
mem['h00EE] = 32'h00050793;
mem['h00EF] = 32'h00078413;
mem['h00F0] = 32'h00812783;
mem['h00F1] = 32'h01878793;
mem['h00F2] = 32'h00078593;
mem['h00F3] = 32'h00040513;
mem['h00F4] = 32'hEA9FF0EF;
mem['h00F5] = 32'h00C12783;
mem['h00F6] = 32'h0087AC23;
mem['h00F7] = 32'h00000013;
mem['h00F8] = 32'h01C12083;
mem['h00F9] = 32'h01812403;
mem['h00FA] = 32'h02010113;
mem['h00FB] = 32'h00008067;
mem['h00FC] = 32'hFF010113;
mem['h00FD] = 32'h00A12623;
mem['h00FE] = 32'h00B12423;
mem['h00FF] = 32'h00C12783;
mem['h0100] = 32'h00812703;
mem['h0101] = 32'h00E7A023;
mem['h0102] = 32'h00000013;
mem['h0103] = 32'h01010113;
mem['h0104] = 32'h00008067;
mem['h0105] = 32'hFF010113;
mem['h0106] = 32'h00A12623;
mem['h0107] = 32'h00B12423;
mem['h0108] = 32'h00C12783;
mem['h0109] = 32'h00812703;
mem['h010A] = 32'h00E7A023;
mem['h010B] = 32'h00000013;
mem['h010C] = 32'h01010113;
mem['h010D] = 32'h00008067;
mem['h010E] = 32'hFF010113;
mem['h010F] = 32'h00A12623;
mem['h0110] = 32'h00B12423;
mem['h0111] = 32'h00C12783;
mem['h0112] = 32'h00812703;
mem['h0113] = 32'h00E7A023;
mem['h0114] = 32'h00000013;
mem['h0115] = 32'h01010113;
mem['h0116] = 32'h00008067;
mem['h0117] = 32'hFF010113;
mem['h0118] = 32'h00A12623;
mem['h0119] = 32'h00B12423;
mem['h011A] = 32'h00C12783;
mem['h011B] = 32'h00812703;
mem['h011C] = 32'h00E7A023;
mem['h011D] = 32'h00000013;
mem['h011E] = 32'h01010113;
mem['h011F] = 32'h00008067;
mem['h0120] = 32'hFF010113;
mem['h0121] = 32'h00A12623;
mem['h0122] = 32'h00B12423;
mem['h0123] = 32'h00C12783;
mem['h0124] = 32'h00812703;
mem['h0125] = 32'h00E7A023;
mem['h0126] = 32'h00000013;
mem['h0127] = 32'h01010113;
mem['h0128] = 32'h00008067;
mem['h0129] = 32'hFF010113;
mem['h012A] = 32'h00A12623;
mem['h012B] = 32'h00B12423;
mem['h012C] = 32'h00C12783;
mem['h012D] = 32'h00812703;
mem['h012E] = 32'h00E7A023;
mem['h012F] = 32'h00000013;
mem['h0130] = 32'h01010113;
mem['h0131] = 32'h00008067;
mem['h0132] = 32'hFF010113;
mem['h0133] = 32'h00A12623;
mem['h0134] = 32'h00B12423;
mem['h0135] = 32'h00C12783;
mem['h0136] = 32'h00812703;
mem['h0137] = 32'h00E7A023;
mem['h0138] = 32'h00000013;
mem['h0139] = 32'h01010113;
mem['h013A] = 32'h00008067;
mem['h013B] = 32'hFE010113;
mem['h013C] = 32'h00112E23;
mem['h013D] = 32'h00812C23;
mem['h013E] = 32'h00A12623;
mem['h013F] = 32'h00B12423;
mem['h0140] = 32'h00400513;
mem['h0141] = 32'hBC1FF0EF;
mem['h0142] = 32'h00050793;
mem['h0143] = 32'h00078413;
mem['h0144] = 32'h00812583;
mem['h0145] = 32'h00040513;
mem['h0146] = 32'hED9FF0EF;
mem['h0147] = 32'h00C12783;
mem['h0148] = 32'h0087A023;
mem['h0149] = 32'h00400513;
mem['h014A] = 32'hB9DFF0EF;
mem['h014B] = 32'h00050793;
mem['h014C] = 32'h00078413;
mem['h014D] = 32'h00812783;
mem['h014E] = 32'h00478793;
mem['h014F] = 32'h00078593;
mem['h0150] = 32'h00040513;
mem['h0151] = 32'hED1FF0EF;
mem['h0152] = 32'h00C12783;
mem['h0153] = 32'h0087A223;
mem['h0154] = 32'h00400513;
mem['h0155] = 32'hB71FF0EF;
mem['h0156] = 32'h00050793;
mem['h0157] = 32'h00078413;
mem['h0158] = 32'h00812783;
mem['h0159] = 32'h00878793;
mem['h015A] = 32'h00078593;
mem['h015B] = 32'h00040513;
mem['h015C] = 32'hEC9FF0EF;
mem['h015D] = 32'h00C12783;
mem['h015E] = 32'h0087A423;
mem['h015F] = 32'h00400513;
mem['h0160] = 32'hB45FF0EF;
mem['h0161] = 32'h00050793;
mem['h0162] = 32'h00078413;
mem['h0163] = 32'h00812783;
mem['h0164] = 32'h00C78793;
mem['h0165] = 32'h00078593;
mem['h0166] = 32'h00040513;
mem['h0167] = 32'hEC1FF0EF;
mem['h0168] = 32'h00C12783;
mem['h0169] = 32'h0087A623;
mem['h016A] = 32'h00400513;
mem['h016B] = 32'hB19FF0EF;
mem['h016C] = 32'h00050793;
mem['h016D] = 32'h00078413;
mem['h016E] = 32'h00812783;
mem['h016F] = 32'h01078793;
mem['h0170] = 32'h00078593;
mem['h0171] = 32'h00040513;
mem['h0172] = 32'hEB9FF0EF;
mem['h0173] = 32'h00C12783;
mem['h0174] = 32'h0087A823;
mem['h0175] = 32'h00400513;
mem['h0176] = 32'hAEDFF0EF;
mem['h0177] = 32'h00050793;
mem['h0178] = 32'h00078413;
mem['h0179] = 32'h00812783;
mem['h017A] = 32'h01478793;
mem['h017B] = 32'h00078593;
mem['h017C] = 32'h00040513;
mem['h017D] = 32'hEB1FF0EF;
mem['h017E] = 32'h00C12783;
mem['h017F] = 32'h0087AA23;
mem['h0180] = 32'h00400513;
mem['h0181] = 32'hAC1FF0EF;
mem['h0182] = 32'h00050793;
mem['h0183] = 32'h00078413;
mem['h0184] = 32'h00812783;
mem['h0185] = 32'h01878793;
mem['h0186] = 32'h00078593;
mem['h0187] = 32'h00040513;
mem['h0188] = 32'hEA9FF0EF;
mem['h0189] = 32'h00C12783;
mem['h018A] = 32'h0087AC23;
mem['h018B] = 32'h00000013;
mem['h018C] = 32'h01C12083;
mem['h018D] = 32'h01812403;
mem['h018E] = 32'h02010113;
mem['h018F] = 32'h00008067;
mem['h0190] = 32'hFE010113;
mem['h0191] = 32'h00112E23;
mem['h0192] = 32'h00812C23;
mem['h0193] = 32'h00A12623;
mem['h0194] = 32'h00B12423;
mem['h0195] = 32'h01C00513;
mem['h0196] = 32'hA6DFF0EF;
mem['h0197] = 32'h00050793;
mem['h0198] = 32'h00078413;
mem['h0199] = 32'h00812583;
mem['h019A] = 32'h00040513;
mem['h019B] = 32'hC31FF0EF;
mem['h019C] = 32'h00C12783;
mem['h019D] = 32'h0087A023;
mem['h019E] = 32'h01C00513;
mem['h019F] = 32'hA49FF0EF;
mem['h01A0] = 32'h00050793;
mem['h01A1] = 32'h00078413;
mem['h01A2] = 32'h00812783;
mem['h01A3] = 32'h01C78793;
mem['h01A4] = 32'h00078593;
mem['h01A5] = 32'h00040513;
mem['h01A6] = 32'hE55FF0EF;
mem['h01A7] = 32'h00C12783;
mem['h01A8] = 32'h0087A223;
mem['h01A9] = 32'h00000013;
mem['h01AA] = 32'h01C12083;
mem['h01AB] = 32'h01812403;
mem['h01AC] = 32'h02010113;
mem['h01AD] = 32'h00008067;
mem['h01AE] = 32'hFF010113;
mem['h01AF] = 32'h00A12623;
mem['h01B0] = 32'h00B12423;
mem['h01B1] = 32'h00C12783;
mem['h01B2] = 32'h00812703;
mem['h01B3] = 32'h00E7A023;
mem['h01B4] = 32'h00000013;
mem['h01B5] = 32'h01010113;
mem['h01B6] = 32'h00008067;
mem['h01B7] = 32'hFF010113;
mem['h01B8] = 32'h00A12623;
mem['h01B9] = 32'h00B12423;
mem['h01BA] = 32'h00C12783;
mem['h01BB] = 32'h00812703;
mem['h01BC] = 32'h00E7A023;
mem['h01BD] = 32'h00000013;
mem['h01BE] = 32'h01010113;
mem['h01BF] = 32'h00008067;
mem['h01C0] = 32'hFF010113;
mem['h01C1] = 32'h00A12623;
mem['h01C2] = 32'h00B12423;
mem['h01C3] = 32'h00C12783;
mem['h01C4] = 32'h00812703;
mem['h01C5] = 32'h00E7A023;
mem['h01C6] = 32'h00000013;
mem['h01C7] = 32'h01010113;
mem['h01C8] = 32'h00008067;
mem['h01C9] = 32'hFF010113;
mem['h01CA] = 32'h00A12623;
mem['h01CB] = 32'h00B12423;
mem['h01CC] = 32'h00C12783;
mem['h01CD] = 32'h00812703;
mem['h01CE] = 32'h00E7A023;
mem['h01CF] = 32'h00000013;
mem['h01D0] = 32'h01010113;
mem['h01D1] = 32'h00008067;
mem['h01D2] = 32'hFE010113;
mem['h01D3] = 32'h00112E23;
mem['h01D4] = 32'h00812C23;
mem['h01D5] = 32'h00A12623;
mem['h01D6] = 32'h00B12423;
mem['h01D7] = 32'h00400513;
mem['h01D8] = 32'h965FF0EF;
mem['h01D9] = 32'h00050793;
mem['h01DA] = 32'h00078413;
mem['h01DB] = 32'h00812583;
mem['h01DC] = 32'h00040513;
mem['h01DD] = 32'hF45FF0EF;
mem['h01DE] = 32'h00C12783;
mem['h01DF] = 32'h0087A023;
mem['h01E0] = 32'h00400513;
mem['h01E1] = 32'h941FF0EF;
mem['h01E2] = 32'h00050793;
mem['h01E3] = 32'h00078413;
mem['h01E4] = 32'h00812783;
mem['h01E5] = 32'h00478793;
mem['h01E6] = 32'h00078593;
mem['h01E7] = 32'h00040513;
mem['h01E8] = 32'hF3DFF0EF;
mem['h01E9] = 32'h00C12783;
mem['h01EA] = 32'h0087A223;
mem['h01EB] = 32'h00400513;
mem['h01EC] = 32'h915FF0EF;
mem['h01ED] = 32'h00050793;
mem['h01EE] = 32'h00078413;
mem['h01EF] = 32'h00812783;
mem['h01F0] = 32'h00878793;
mem['h01F1] = 32'h00078593;
mem['h01F2] = 32'h00040513;
mem['h01F3] = 32'hF35FF0EF;
mem['h01F4] = 32'h00C12783;
mem['h01F5] = 32'h0087A423;
mem['h01F6] = 32'h00400513;
mem['h01F7] = 32'h8E9FF0EF;
mem['h01F8] = 32'h00050793;
mem['h01F9] = 32'h00078413;
mem['h01FA] = 32'h00812783;
mem['h01FB] = 32'h00C78793;
mem['h01FC] = 32'h00078593;
mem['h01FD] = 32'h00040513;
mem['h01FE] = 32'hF2DFF0EF;
mem['h01FF] = 32'h00C12783;
mem['h0200] = 32'h0087A623;
mem['h0201] = 32'h00000013;
mem['h0202] = 32'h01C12083;
mem['h0203] = 32'h01812403;
mem['h0204] = 32'h02010113;
mem['h0205] = 32'h00008067;
mem['h0206] = 32'hFF010113;
mem['h0207] = 32'h00A12623;
mem['h0208] = 32'h00B12423;
mem['h0209] = 32'h00C12783;
mem['h020A] = 32'h00812703;
mem['h020B] = 32'h00E7A023;
mem['h020C] = 32'h00000013;
mem['h020D] = 32'h01010113;
mem['h020E] = 32'h00008067;
mem['h020F] = 32'hFF010113;
mem['h0210] = 32'h00A12623;
mem['h0211] = 32'h00B12423;
mem['h0212] = 32'h00C12783;
mem['h0213] = 32'h00812703;
mem['h0214] = 32'h00E7A023;
mem['h0215] = 32'h00000013;
mem['h0216] = 32'h01010113;
mem['h0217] = 32'h00008067;
mem['h0218] = 32'hFE010113;
mem['h0219] = 32'h00112E23;
mem['h021A] = 32'h00812C23;
mem['h021B] = 32'h00A12623;
mem['h021C] = 32'h00B12423;
mem['h021D] = 32'h00400513;
mem['h021E] = 32'h84DFF0EF;
mem['h021F] = 32'h00050793;
mem['h0220] = 32'h00078413;
mem['h0221] = 32'h00812583;
mem['h0222] = 32'h00040513;
mem['h0223] = 32'hFB1FF0EF;
mem['h0224] = 32'h00C12783;
mem['h0225] = 32'h0087A023;
mem['h0226] = 32'h00000013;
mem['h0227] = 32'h01C12083;
mem['h0228] = 32'h01812403;
mem['h0229] = 32'h02010113;
mem['h022A] = 32'h00008067;
mem['h022B] = 32'hFF010113;
mem['h022C] = 32'h00A12623;
mem['h022D] = 32'h00B12423;
mem['h022E] = 32'h00C12783;
mem['h022F] = 32'h00812703;
mem['h0230] = 32'h00E7A023;
mem['h0231] = 32'h00000013;
mem['h0232] = 32'h01010113;
mem['h0233] = 32'h00008067;
mem['h0234] = 32'hFE010113;
mem['h0235] = 32'h00112E23;
mem['h0236] = 32'h00812C23;
mem['h0237] = 32'h00A12623;
mem['h0238] = 32'h00B12423;
mem['h0239] = 32'h00400513;
mem['h023A] = 32'hFDCFF0EF;
mem['h023B] = 32'h00050793;
mem['h023C] = 32'h00078413;
mem['h023D] = 32'h00812583;
mem['h023E] = 32'h00040513;
mem['h023F] = 32'hFB1FF0EF;
mem['h0240] = 32'h00C12783;
mem['h0241] = 32'h0087A023;
mem['h0242] = 32'h00000013;
mem['h0243] = 32'h01C12083;
mem['h0244] = 32'h01812403;
mem['h0245] = 32'h02010113;
mem['h0246] = 32'h00008067;
mem['h0247] = 32'hFF010113;
mem['h0248] = 32'h00A12623;
mem['h0249] = 32'h00B12423;
mem['h024A] = 32'h00C12783;
mem['h024B] = 32'h00812703;
mem['h024C] = 32'h00E7A023;
mem['h024D] = 32'h00000013;
mem['h024E] = 32'h01010113;
mem['h024F] = 32'h00008067;
mem['h0250] = 32'hFD010113;
mem['h0251] = 32'h02112623;
mem['h0252] = 32'h02812423;
mem['h0253] = 32'h00A12623;
mem['h0254] = 32'h00B12423;
mem['h0255] = 32'h00800513;
mem['h0256] = 32'hF6CFF0EF;
mem['h0257] = 32'h00050793;
mem['h0258] = 32'h00078413;
mem['h0259] = 32'h00812583;
mem['h025A] = 32'h00040513;
mem['h025B] = 32'hCD5FF0EF;
mem['h025C] = 32'h00C12783;
mem['h025D] = 32'h0087A023;
mem['h025E] = 32'h01000513;
mem['h025F] = 32'hF48FF0EF;
mem['h0260] = 32'h00050793;
mem['h0261] = 32'h00078413;
mem['h0262] = 32'h00812783;
mem['h0263] = 32'h03878793;
mem['h0264] = 32'h00078593;
mem['h0265] = 32'h00040513;
mem['h0266] = 32'hDB1FF0EF;
mem['h0267] = 32'h00C12783;
mem['h0268] = 32'h0087A223;
mem['h0269] = 32'h00400513;
mem['h026A] = 32'hF1CFF0EF;
mem['h026B] = 32'h00050793;
mem['h026C] = 32'h00078413;
mem['h026D] = 32'h00812783;
mem['h026E] = 32'h04878793;
mem['h026F] = 32'h00078593;
mem['h0270] = 32'h00040513;
mem['h0271] = 32'hE55FF0EF;
mem['h0272] = 32'h00C12783;
mem['h0273] = 32'h0087A423;
mem['h0274] = 32'h00012E23;
mem['h0275] = 32'h0540006F;
mem['h0276] = 32'h00400513;
mem['h0277] = 32'hEE8FF0EF;
mem['h0278] = 32'h00050793;
mem['h0279] = 32'h00078413;
mem['h027A] = 32'h01C12783;
mem['h027B] = 32'h01378793;
mem['h027C] = 32'h00279793;
mem['h027D] = 32'h00812703;
mem['h027E] = 32'h00F707B3;
mem['h027F] = 32'h00078593;
mem['h0280] = 32'h00040513;
mem['h0281] = 32'hE5DFF0EF;
mem['h0282] = 32'h00C12703;
mem['h0283] = 32'h01C12783;
mem['h0284] = 32'h00279793;
mem['h0285] = 32'h00F707B3;
mem['h0286] = 32'h0087A623;
mem['h0287] = 32'h01C12783;
mem['h0288] = 32'h00178793;
mem['h0289] = 32'h00F12E23;
mem['h028A] = 32'h01C12703;
mem['h028B] = 32'h00300793;
mem['h028C] = 32'hFAE7D4E3;
mem['h028D] = 32'h00400513;
mem['h028E] = 32'hE8CFF0EF;
mem['h028F] = 32'h00050793;
mem['h0290] = 32'h00078413;
mem['h0291] = 32'h00812783;
mem['h0292] = 32'h05C78793;
mem['h0293] = 32'h00078593;
mem['h0294] = 32'h00040513;
mem['h0295] = 32'hE7DFF0EF;
mem['h0296] = 32'h00C12783;
mem['h0297] = 32'h0087AE23;
mem['h0298] = 32'h00400513;
mem['h0299] = 32'hE60FF0EF;
mem['h029A] = 32'h00050793;
mem['h029B] = 32'h00078413;
mem['h029C] = 32'h00812783;
mem['h029D] = 32'h06078793;
mem['h029E] = 32'h00078593;
mem['h029F] = 32'h00040513;
mem['h02A0] = 32'hE9DFF0EF;
mem['h02A1] = 32'h00C12783;
mem['h02A2] = 32'h0287A023;
mem['h02A3] = 32'h00000013;
mem['h02A4] = 32'h02C12083;
mem['h02A5] = 32'h02812403;
mem['h02A6] = 32'h03010113;
mem['h02A7] = 32'h00008067;
mem['h02A8] = 32'hFE010113;
mem['h02A9] = 32'h00112E23;
mem['h02AA] = 32'h00A12623;
mem['h02AB] = 32'h00058793;
mem['h02AC] = 32'h00F105A3;
mem['h02AD] = 32'h00000013;
mem['h02AE] = 32'h00C12783;
mem['h02AF] = 32'h0047A783;
mem['h02B0] = 32'h0087A783;
mem['h02B1] = 32'h00078513;
mem['h02B2] = 32'h388000EF;
mem['h02B3] = 32'h00050793;
mem['h02B4] = 32'h00F037B3;
mem['h02B5] = 32'h0FF7F793;
mem['h02B6] = 32'hFE0790E3;
mem['h02B7] = 32'h00C12783;
mem['h02B8] = 32'h0047A783;
mem['h02B9] = 32'h0087A783;
mem['h02BA] = 32'h00B14703;
mem['h02BB] = 32'h00070593;
mem['h02BC] = 32'h00078513;
mem['h02BD] = 32'h330000EF;
mem['h02BE] = 32'h00000013;
mem['h02BF] = 32'h01C12083;
mem['h02C0] = 32'h02010113;
mem['h02C1] = 32'h00008067;
mem['h02C2] = 32'hFD010113;
mem['h02C3] = 32'h02112623;
mem['h02C4] = 32'h00A12623;
mem['h02C5] = 32'h00B12423;
mem['h02C6] = 32'h00C12223;
mem['h02C7] = 32'h00412783;
mem['h02C8] = 32'hFFF78793;
mem['h02C9] = 32'h00279793;
mem['h02CA] = 32'h00F12E23;
mem['h02CB] = 32'h03C0006F;
mem['h02CC] = 32'h01C12783;
mem['h02CD] = 32'h00812703;
mem['h02CE] = 32'h00F757B3;
mem['h02CF] = 32'h00F7F793;
mem['h02D0] = 32'h00001737;
mem['h02D1] = 32'h07C70713;
mem['h02D2] = 32'h00F707B3;
mem['h02D3] = 32'h0007C783;
mem['h02D4] = 32'h00078593;
mem['h02D5] = 32'h00C12503;
mem['h02D6] = 32'hF49FF0EF;
mem['h02D7] = 32'h01C12783;
mem['h02D8] = 32'hFFC78793;
mem['h02D9] = 32'h00F12E23;
mem['h02DA] = 32'h01C12783;
mem['h02DB] = 32'hFC07D2E3;
mem['h02DC] = 32'h00000013;
mem['h02DD] = 32'h00000013;
mem['h02DE] = 32'h02C12083;
mem['h02DF] = 32'h03010113;
mem['h02E0] = 32'h00008067;
mem['h02E1] = 32'hFE010113;
mem['h02E2] = 32'h00112E23;
mem['h02E3] = 32'h00A12623;
mem['h02E4] = 32'h00B12423;
mem['h02E5] = 32'h0200006F;
mem['h02E6] = 32'h00812783;
mem['h02E7] = 32'h00178713;
mem['h02E8] = 32'h00E12423;
mem['h02E9] = 32'h0007C783;
mem['h02EA] = 32'h00078593;
mem['h02EB] = 32'h00C12503;
mem['h02EC] = 32'hEF1FF0EF;
mem['h02ED] = 32'h00812783;
mem['h02EE] = 32'h0007C783;
mem['h02EF] = 32'hFC079EE3;
mem['h02F0] = 32'h00000013;
mem['h02F1] = 32'h00000013;
mem['h02F2] = 32'h01C12083;
mem['h02F3] = 32'h02010113;
mem['h02F4] = 32'h00008067;
mem['h02F5] = 32'hFD010113;
mem['h02F6] = 32'h02112623;
mem['h02F7] = 32'h00A12623;
mem['h02F8] = 32'h00B12423;
mem['h02F9] = 32'h00012E23;
mem['h02FA] = 32'h0D00006F;
mem['h02FB] = 32'h00C12783;
mem['h02FC] = 32'h0047A783;
mem['h02FD] = 32'h0007A783;
mem['h02FE] = 32'h00078513;
mem['h02FF] = 32'h208000EF;
mem['h0300] = 32'h00A12C23;
mem['h0301] = 32'h01812783;
mem['h0302] = 32'hFE07D2E3;
mem['h0303] = 32'h01812783;
mem['h0304] = 32'h0FF7F713;
mem['h0305] = 32'h00812783;
mem['h0306] = 32'h00E78023;
mem['h0307] = 32'h00812783;
mem['h0308] = 32'h0007C783;
mem['h0309] = 32'h00078593;
mem['h030A] = 32'h00C12503;
mem['h030B] = 32'hE75FF0EF;
mem['h030C] = 32'h01C12703;
mem['h030D] = 32'h01D00793;
mem['h030E] = 32'h04F71063;
mem['h030F] = 32'h00812783;
mem['h0310] = 32'h00D00713;
mem['h0311] = 32'h00E78023;
mem['h0312] = 32'h00812783;
mem['h0313] = 32'h00178793;
mem['h0314] = 32'h00F12423;
mem['h0315] = 32'h00812783;
mem['h0316] = 32'h00A00713;
mem['h0317] = 32'h00E78023;
mem['h0318] = 32'h00812783;
mem['h0319] = 32'h00178793;
mem['h031A] = 32'h00F12423;
mem['h031B] = 32'h00812783;
mem['h031C] = 32'h00078023;
mem['h031D] = 32'h0540006F;
mem['h031E] = 32'h00812783;
mem['h031F] = 32'h0007C703;
mem['h0320] = 32'h00A00793;
mem['h0321] = 32'h00F71E63;
mem['h0322] = 32'h00812783;
mem['h0323] = 32'h00178793;
mem['h0324] = 32'h00F12423;
mem['h0325] = 32'h00812783;
mem['h0326] = 32'h00078023;
mem['h0327] = 32'h02C0006F;
mem['h0328] = 32'h00812783;
mem['h0329] = 32'h00178793;
mem['h032A] = 32'h00F12423;
mem['h032B] = 32'h01C12783;
mem['h032C] = 32'h00178793;
mem['h032D] = 32'h00F12E23;
mem['h032E] = 32'h01C12703;
mem['h032F] = 32'h01E00793;
mem['h0330] = 32'hF2E7D6E3;
mem['h0331] = 32'h00000013;
mem['h0332] = 32'h00000013;
mem['h0333] = 32'h02C12083;
mem['h0334] = 32'h03010113;
mem['h0335] = 32'h00008067;
mem['h0336] = 32'hFB010113;
mem['h0337] = 32'h04112623;
mem['h0338] = 32'h00A12623;
mem['h0339] = 32'h000017B7;
mem['h033A] = 32'h09078793;
mem['h033B] = 32'h02F12C23;
mem['h033C] = 32'h000017B7;
mem['h033D] = 32'h0A478593;
mem['h033E] = 32'h00C12503;
mem['h033F] = 32'hE89FF0EF;
mem['h0340] = 32'h000017B7;
mem['h0341] = 32'h0C078593;
mem['h0342] = 32'h00C12503;
mem['h0343] = 32'hE79FF0EF;
mem['h0344] = 32'h00300793;
mem['h0345] = 32'h02F12E23;
mem['h0346] = 32'h0C40006F;
mem['h0347] = 32'h01410793;
mem['h0348] = 32'h02F12A23;
mem['h0349] = 32'h03412583;
mem['h034A] = 32'h00C12503;
mem['h034B] = 32'hEA9FF0EF;
mem['h034C] = 32'h000017B7;
mem['h034D] = 32'h10078593;
mem['h034E] = 32'h00C12503;
mem['h034F] = 32'hE49FF0EF;
mem['h0350] = 32'h03412583;
mem['h0351] = 32'h00C12503;
mem['h0352] = 32'hE3DFF0EF;
mem['h0353] = 32'h03412583;
mem['h0354] = 32'h03812503;
mem['h0355] = 32'h2D8000EF;
mem['h0356] = 32'h00050793;
mem['h0357] = 32'h0017B793;
mem['h0358] = 32'h0FF7F793;
mem['h0359] = 32'h00078C63;
mem['h035A] = 32'h000017B7;
mem['h035B] = 32'h11478593;
mem['h035C] = 32'h00C12503;
mem['h035D] = 32'hE11FF0EF;
mem['h035E] = 32'h06C0006F;
mem['h035F] = 32'h000017B7;
mem['h0360] = 32'h12C78593;
mem['h0361] = 32'h00C12503;
mem['h0362] = 32'hDFDFF0EF;
mem['h0363] = 32'h03C12703;
mem['h0364] = 32'h00100793;
mem['h0365] = 32'h02E7DE63;
mem['h0366] = 32'h000017B7;
mem['h0367] = 32'h14878593;
mem['h0368] = 32'h00C12503;
mem['h0369] = 32'hDE1FF0EF;
mem['h036A] = 32'h03C12783;
mem['h036B] = 32'hFFF78793;
mem['h036C] = 32'h00100613;
mem['h036D] = 32'h00078593;
mem['h036E] = 32'h00C12503;
mem['h036F] = 32'hD4DFF0EF;
mem['h0370] = 32'h000017B7;
mem['h0371] = 32'h16C78593;
mem['h0372] = 32'h00C12503;
mem['h0373] = 32'hDB9FF0EF;
mem['h0374] = 32'h03C12783;
mem['h0375] = 32'hFFF78793;
mem['h0376] = 32'h02F12E23;
mem['h0377] = 32'h03C12783;
mem['h0378] = 32'hF2F04EE3;
mem['h0379] = 32'h000017B7;
mem['h037A] = 32'h17478593;
mem['h037B] = 32'h00C12503;
mem['h037C] = 32'hD95FF0EF;
mem['h037D] = 32'h00000013;
mem['h037E] = 32'h04C12083;
mem['h037F] = 32'h05010113;
mem['h0380] = 32'h00008067;
mem['h0381] = 32'hFF010113;
mem['h0382] = 32'h00A12623;
mem['h0383] = 32'h00C12783;
mem['h0384] = 32'h0007A783;
mem['h0385] = 32'h0007A783;
mem['h0386] = 32'h00078513;
mem['h0387] = 32'h01010113;
mem['h0388] = 32'h00008067;
mem['h0389] = 32'hFF010113;
mem['h038A] = 32'h00A12623;
mem['h038B] = 32'h00B12423;
mem['h038C] = 32'h00C12783;
mem['h038D] = 32'h0007A783;
mem['h038E] = 32'h00812703;
mem['h038F] = 32'h0FF77713;
mem['h0390] = 32'h00E78023;
mem['h0391] = 32'h00000013;
mem['h0392] = 32'h01010113;
mem['h0393] = 32'h00008067;
mem['h0394] = 32'hFF010113;
mem['h0395] = 32'h00A12623;
mem['h0396] = 32'h00C12783;
mem['h0397] = 32'h0007A783;
mem['h0398] = 32'h0007A783;
mem['h0399] = 32'h01F7D793;
mem['h039A] = 32'h0FF7F793;
mem['h039B] = 32'h00078513;
mem['h039C] = 32'h01010113;
mem['h039D] = 32'h00008067;
mem['h039E] = 32'hFE010113;
mem['h039F] = 32'h00A12623;
mem['h03A0] = 32'h00B12423;
mem['h03A1] = 32'h00C12223;
mem['h03A2] = 32'h00C12783;
mem['h03A3] = 32'h00F12C23;
mem['h03A4] = 32'h00812783;
mem['h03A5] = 32'h00F10BA3;
mem['h03A6] = 32'h00012E23;
mem['h03A7] = 32'h0240006F;
mem['h03A8] = 32'h01812703;
mem['h03A9] = 32'h01C12783;
mem['h03AA] = 32'h00F707B3;
mem['h03AB] = 32'h01714703;
mem['h03AC] = 32'h00E78023;
mem['h03AD] = 32'h01C12783;
mem['h03AE] = 32'h00178793;
mem['h03AF] = 32'h00F12E23;
mem['h03B0] = 32'h01C12703;
mem['h03B1] = 32'h00412783;
mem['h03B2] = 32'hFCF76CE3;
mem['h03B3] = 32'h00C12783;
mem['h03B4] = 32'h00078513;
mem['h03B5] = 32'h02010113;
mem['h03B6] = 32'h00008067;
mem['h03B7] = 32'hFE010113;
mem['h03B8] = 32'h00A12623;
mem['h03B9] = 32'h00B12423;
mem['h03BA] = 32'h00C12223;
mem['h03BB] = 32'h00C12783;
mem['h03BC] = 32'h00F12C23;
mem['h03BD] = 32'h00812783;
mem['h03BE] = 32'h00F12A23;
mem['h03BF] = 32'h00012E23;
mem['h03C0] = 32'h0300006F;
mem['h03C1] = 32'h01412703;
mem['h03C2] = 32'h01C12783;
mem['h03C3] = 32'h00F70733;
mem['h03C4] = 32'h01812683;
mem['h03C5] = 32'h01C12783;
mem['h03C6] = 32'h00F687B3;
mem['h03C7] = 32'h00074703;
mem['h03C8] = 32'h00E78023;
mem['h03C9] = 32'h01C12783;
mem['h03CA] = 32'h00178793;
mem['h03CB] = 32'h00F12E23;
mem['h03CC] = 32'h01C12703;
mem['h03CD] = 32'h00412783;
mem['h03CE] = 32'hFCF766E3;
mem['h03CF] = 32'h00C12783;
mem['h03D0] = 32'h00078513;
mem['h03D1] = 32'h02010113;
mem['h03D2] = 32'h00008067;
mem['h03D3] = 32'hFE010113;
mem['h03D4] = 32'h00A12623;
mem['h03D5] = 32'h00B12423;
mem['h03D6] = 32'h00C12223;
mem['h03D7] = 32'h00C12783;
mem['h03D8] = 32'h00F12C23;
mem['h03D9] = 32'h00812783;
mem['h03DA] = 32'h00F12A23;
mem['h03DB] = 32'h00012E23;
mem['h03DC] = 32'h0600006F;
mem['h03DD] = 32'h01812703;
mem['h03DE] = 32'h01C12783;
mem['h03DF] = 32'h00F707B3;
mem['h03E0] = 32'h0007C703;
mem['h03E1] = 32'h01412683;
mem['h03E2] = 32'h01C12783;
mem['h03E3] = 32'h00F687B3;
mem['h03E4] = 32'h0007C783;
mem['h03E5] = 32'h02F70863;
mem['h03E6] = 32'h01812703;
mem['h03E7] = 32'h01C12783;
mem['h03E8] = 32'h00F707B3;
mem['h03E9] = 32'h0007C783;
mem['h03EA] = 32'h00078693;
mem['h03EB] = 32'h01412703;
mem['h03EC] = 32'h01C12783;
mem['h03ED] = 32'h00F707B3;
mem['h03EE] = 32'h0007C783;
mem['h03EF] = 32'h40F687B3;
mem['h03F0] = 32'h0200006F;
mem['h03F1] = 32'h01C12783;
mem['h03F2] = 32'h00178793;
mem['h03F3] = 32'h00F12E23;
mem['h03F4] = 32'h01C12703;
mem['h03F5] = 32'h00412783;
mem['h03F6] = 32'hF8F76EE3;
mem['h03F7] = 32'h00000793;
mem['h03F8] = 32'h00078513;
mem['h03F9] = 32'h02010113;
mem['h03FA] = 32'h00008067;
mem['h03FB] = 32'hFE010113;
mem['h03FC] = 32'h00A12623;
mem['h03FD] = 32'h00012E23;
mem['h03FE] = 32'h0100006F;
mem['h03FF] = 32'h01C12783;
mem['h0400] = 32'h00178793;
mem['h0401] = 32'h00F12E23;
mem['h0402] = 32'h00C12703;
mem['h0403] = 32'h01C12783;
mem['h0404] = 32'h00F707B3;
mem['h0405] = 32'h0007C783;
mem['h0406] = 32'hFE0792E3;
mem['h0407] = 32'h01C12783;
mem['h0408] = 32'h00078513;
mem['h0409] = 32'h02010113;
mem['h040A] = 32'h00008067;
mem['h040B] = 32'hFE010113;
mem['h040C] = 32'h00112E23;
mem['h040D] = 32'h00A12623;
mem['h040E] = 32'h00B12423;
mem['h040F] = 32'h00C12503;
mem['h0410] = 32'hFADFF0EF;
mem['h0411] = 32'h00050793;
mem['h0412] = 32'h00078613;
mem['h0413] = 32'h00812583;
mem['h0414] = 32'h00C12503;
mem['h0415] = 32'hEF9FF0EF;
mem['h0416] = 32'h00050793;
mem['h0417] = 32'h00078513;
mem['h0418] = 32'h01C12083;
mem['h0419] = 32'h02010113;
mem['h041A] = 32'h00008067;
mem['h041B] = 32'h6C6C6548;
mem['h041C] = 32'h6F77206F;
mem['h041D] = 32'h21646C72;
mem['h041E] = 32'h00000A0D;
mem['h041F] = 32'h33323130;
mem['h0420] = 32'h37363534;
mem['h0421] = 32'h42413938;
mem['h0422] = 32'h46454443;
mem['h0423] = 32'h00000000;
mem['h0424] = 32'h7320694D;
mem['h0425] = 32'h46206F6D;
mem['h0426] = 32'h20414750;
mem['h0427] = 32'h616A6172;
mem['h0428] = 32'h00000A0D;
mem['h0429] = 32'h530A0A0D;
mem['h042A] = 32'h6D616C65;
mem['h042B] = 32'h75646520;
mem['h042C] = 32'h20434F53;
mem['h042D] = 32'h6B636148;
mem['h042E] = 32'h21737265;
mem['h042F] = 32'h00000A0D;
mem['h0430] = 32'h20797254;
mem['h0431] = 32'h73657567;
mem['h0432] = 32'h676E6973;
mem['h0433] = 32'h74203320;
mem['h0434] = 32'h73656D69;
mem['h0435] = 32'h61687720;
mem['h0436] = 32'h27492074;
mem['h0437] = 32'h6874206D;
mem['h0438] = 32'h696B6E69;
mem['h0439] = 32'h202C676E;
mem['h043A] = 32'h6E656874;
mem['h043B] = 32'h65727020;
mem['h043C] = 32'h3C207373;
mem['h043D] = 32'h45544E45;
mem['h043E] = 32'h0D2E3E52;
mem['h043F] = 32'h0000000A;
mem['h0440] = 32'h090A0A0D;
mem['h0441] = 32'h20756F59;
mem['h0442] = 32'h65746E65;
mem['h0443] = 32'h3A646572;
mem['h0444] = 32'h00000020;
mem['h0445] = 32'h7C090A0D;
mem['h0446] = 32'h756F5920;
mem['h0447] = 32'h74696820;
mem['h0448] = 32'h21746920;
mem['h0449] = 32'h292D3A20;
mem['h044A] = 32'h00000A0D;
mem['h044B] = 32'h7C090A0D;
mem['h044C] = 32'h726F5320;
mem['h044D] = 32'h202C7972;
mem['h044E] = 32'h20756F79;
mem['h044F] = 32'h7373696D;
mem['h0450] = 32'h69206465;
mem['h0451] = 32'h00002E74;
mem['h0452] = 32'h7C090A0D;
mem['h0453] = 32'h2E2E2E20;
mem['h0454] = 32'h20797254;
mem['h0455] = 32'h69616761;
mem['h0456] = 32'h43202E6E;
mem['h0457] = 32'h69646572;
mem['h0458] = 32'h656C2074;
mem['h0459] = 32'h203A7466;
mem['h045A] = 32'h00000000;
mem['h045B] = 32'h0A0A0A0D;
mem['h045C] = 32'h00000000;
mem['h045D] = 32'h4F440A0D;
mem['h045E] = 32'h0D21454E;
mem['h045F] = 32'h0000000A;
