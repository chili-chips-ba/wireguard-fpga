mem['h0000] = 32'h00002517;
mem['h0001] = 32'h75850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h60C18593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h420020EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'hFF010113;
mem['h001D] = 32'h00A12623;
mem['h001E] = 32'h00C12783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'h0007A783;
mem['h0021] = 32'h00078513;
mem['h0022] = 32'h01010113;
mem['h0023] = 32'h00008067;
mem['h0024] = 32'hFF010113;
mem['h0025] = 32'h00A12623;
mem['h0026] = 32'h00B12423;
mem['h0027] = 32'h00C12783;
mem['h0028] = 32'h0007A783;
mem['h0029] = 32'h00812703;
mem['h002A] = 32'h0FF77713;
mem['h002B] = 32'h00E78023;
mem['h002C] = 32'h00000013;
mem['h002D] = 32'h01010113;
mem['h002E] = 32'h00008067;
mem['h002F] = 32'hFF010113;
mem['h0030] = 32'h00A12623;
mem['h0031] = 32'h00C12783;
mem['h0032] = 32'h0007A783;
mem['h0033] = 32'h0007A783;
mem['h0034] = 32'h01F7D793;
mem['h0035] = 32'h0FF7F793;
mem['h0036] = 32'h00078513;
mem['h0037] = 32'h01010113;
mem['h0038] = 32'h00008067;
mem['h0039] = 32'hFE010113;
mem['h003A] = 32'h00112E23;
mem['h003B] = 32'h00A12623;
mem['h003C] = 32'h00058793;
mem['h003D] = 32'h00F105A3;
mem['h003E] = 32'h00000013;
mem['h003F] = 32'h00C12783;
mem['h0040] = 32'h0047A783;
mem['h0041] = 32'h0087A783;
mem['h0042] = 32'h00078513;
mem['h0043] = 32'hFB1FF0EF;
mem['h0044] = 32'h00050793;
mem['h0045] = 32'h00F037B3;
mem['h0046] = 32'h0FF7F793;
mem['h0047] = 32'hFE0790E3;
mem['h0048] = 32'h00C12783;
mem['h0049] = 32'h0047A783;
mem['h004A] = 32'h0087A783;
mem['h004B] = 32'h00B14703;
mem['h004C] = 32'h00070593;
mem['h004D] = 32'h00078513;
mem['h004E] = 32'hF59FF0EF;
mem['h004F] = 32'h00000013;
mem['h0050] = 32'h01C12083;
mem['h0051] = 32'h02010113;
mem['h0052] = 32'h00008067;
mem['h0053] = 32'hFD010113;
mem['h0054] = 32'h02112623;
mem['h0055] = 32'h00A12623;
mem['h0056] = 32'h00B12423;
mem['h0057] = 32'h00C12223;
mem['h0058] = 32'h00412783;
mem['h0059] = 32'hFFF78793;
mem['h005A] = 32'h00279793;
mem['h005B] = 32'h00F12E23;
mem['h005C] = 32'h03C0006F;
mem['h005D] = 32'h01C12783;
mem['h005E] = 32'h00812703;
mem['h005F] = 32'h00F757B3;
mem['h0060] = 32'h00F7F793;
mem['h0061] = 32'h00002737;
mem['h0062] = 32'h64470713;
mem['h0063] = 32'h00F707B3;
mem['h0064] = 32'h0007C783;
mem['h0065] = 32'h00078593;
mem['h0066] = 32'h00C12503;
mem['h0067] = 32'hF49FF0EF;
mem['h0068] = 32'h01C12783;
mem['h0069] = 32'hFFC78793;
mem['h006A] = 32'h00F12E23;
mem['h006B] = 32'h01C12783;
mem['h006C] = 32'hFC07D2E3;
mem['h006D] = 32'h00000013;
mem['h006E] = 32'h00000013;
mem['h006F] = 32'h02C12083;
mem['h0070] = 32'h03010113;
mem['h0071] = 32'h00008067;
mem['h0072] = 32'hFD010113;
mem['h0073] = 32'h02112623;
mem['h0074] = 32'h00A12623;
mem['h0075] = 32'h00058793;
mem['h0076] = 32'h00F11523;
mem['h0077] = 32'h00A15783;
mem['h0078] = 32'h00079A63;
mem['h0079] = 32'h03000593;
mem['h007A] = 32'h00C12503;
mem['h007B] = 32'hEF9FF0EF;
mem['h007C] = 32'h0DC0006F;
mem['h007D] = 32'h00100793;
mem['h007E] = 32'h00F11F23;
mem['h007F] = 32'h0200006F;
mem['h0080] = 32'h01E15783;
mem['h0081] = 32'h00078713;
mem['h0082] = 32'h00070793;
mem['h0083] = 32'h00279793;
mem['h0084] = 32'h00E787B3;
mem['h0085] = 32'h00179793;
mem['h0086] = 32'h00F11F23;
mem['h0087] = 32'h00A15783;
mem['h0088] = 32'h00A00593;
mem['h0089] = 32'h00078513;
mem['h008A] = 32'h370020EF;
mem['h008B] = 32'h00050793;
mem['h008C] = 32'h01079793;
mem['h008D] = 32'h0107D793;
mem['h008E] = 32'h01E15703;
mem['h008F] = 32'hFCE7F2E3;
mem['h0090] = 32'h0840006F;
mem['h0091] = 32'h00A15783;
mem['h0092] = 32'h01E15703;
mem['h0093] = 32'h00070593;
mem['h0094] = 32'h00078513;
mem['h0095] = 32'h344020EF;
mem['h0096] = 32'h00050793;
mem['h0097] = 32'h00F11E23;
mem['h0098] = 32'h01C15783;
mem['h0099] = 32'h0FF7F793;
mem['h009A] = 32'h03078793;
mem['h009B] = 32'h0FF7F793;
mem['h009C] = 32'h00078593;
mem['h009D] = 32'h00C12503;
mem['h009E] = 32'hE6DFF0EF;
mem['h009F] = 32'h01C15783;
mem['h00A0] = 32'h00078713;
mem['h00A1] = 32'h01E15783;
mem['h00A2] = 32'h00078593;
mem['h00A3] = 32'h00070513;
mem['h00A4] = 32'h2DC020EF;
mem['h00A5] = 32'h00050793;
mem['h00A6] = 32'h01079793;
mem['h00A7] = 32'h0107D793;
mem['h00A8] = 32'h00A15703;
mem['h00A9] = 32'h40F707B3;
mem['h00AA] = 32'h00F11523;
mem['h00AB] = 32'h01E15783;
mem['h00AC] = 32'h00A00593;
mem['h00AD] = 32'h00078513;
mem['h00AE] = 32'h2E0020EF;
mem['h00AF] = 32'h00050793;
mem['h00B0] = 32'h00F11F23;
mem['h00B1] = 32'h01E15783;
mem['h00B2] = 32'hF6079EE3;
mem['h00B3] = 32'h02C12083;
mem['h00B4] = 32'h03010113;
mem['h00B5] = 32'h00008067;
mem['h00B6] = 32'hFE010113;
mem['h00B7] = 32'h00112E23;
mem['h00B8] = 32'h00A12623;
mem['h00B9] = 32'h00B12423;
mem['h00BA] = 32'h0200006F;
mem['h00BB] = 32'h00812783;
mem['h00BC] = 32'h00178713;
mem['h00BD] = 32'h00E12423;
mem['h00BE] = 32'h0007C783;
mem['h00BF] = 32'h00078593;
mem['h00C0] = 32'h00C12503;
mem['h00C1] = 32'hDE1FF0EF;
mem['h00C2] = 32'h00812783;
mem['h00C3] = 32'h0007C783;
mem['h00C4] = 32'hFC079EE3;
mem['h00C5] = 32'h00000013;
mem['h00C6] = 32'h00000013;
mem['h00C7] = 32'h01C12083;
mem['h00C8] = 32'h02010113;
mem['h00C9] = 32'h00008067;
mem['h00CA] = 32'hFE010113;
mem['h00CB] = 32'h00112E23;
mem['h00CC] = 32'h00A12623;
mem['h00CD] = 32'h00B12423;
mem['h00CE] = 32'h00812783;
mem['h00CF] = 32'h0007C783;
mem['h00D0] = 32'h00078593;
mem['h00D1] = 32'h00C12503;
mem['h00D2] = 32'hE81FF0EF;
mem['h00D3] = 32'h02E00593;
mem['h00D4] = 32'h00C12503;
mem['h00D5] = 32'hD91FF0EF;
mem['h00D6] = 32'h00812783;
mem['h00D7] = 32'h00178793;
mem['h00D8] = 32'h0007C783;
mem['h00D9] = 32'h00078593;
mem['h00DA] = 32'h00C12503;
mem['h00DB] = 32'hE5DFF0EF;
mem['h00DC] = 32'h02E00593;
mem['h00DD] = 32'h00C12503;
mem['h00DE] = 32'hD6DFF0EF;
mem['h00DF] = 32'h00812783;
mem['h00E0] = 32'h00278793;
mem['h00E1] = 32'h0007C783;
mem['h00E2] = 32'h00078593;
mem['h00E3] = 32'h00C12503;
mem['h00E4] = 32'hE39FF0EF;
mem['h00E5] = 32'h02E00593;
mem['h00E6] = 32'h00C12503;
mem['h00E7] = 32'hD49FF0EF;
mem['h00E8] = 32'h00812783;
mem['h00E9] = 32'h00378793;
mem['h00EA] = 32'h0007C783;
mem['h00EB] = 32'h00078593;
mem['h00EC] = 32'h00C12503;
mem['h00ED] = 32'hE15FF0EF;
mem['h00EE] = 32'h00000013;
mem['h00EF] = 32'h01C12083;
mem['h00F0] = 32'h02010113;
mem['h00F1] = 32'h00008067;
mem['h00F2] = 32'hFE010113;
mem['h00F3] = 32'h00112E23;
mem['h00F4] = 32'h00A12623;
mem['h00F5] = 32'h00B12423;
mem['h00F6] = 32'h00812783;
mem['h00F7] = 32'h0007C783;
mem['h00F8] = 32'h00200613;
mem['h00F9] = 32'h00078593;
mem['h00FA] = 32'h00C12503;
mem['h00FB] = 32'hD61FF0EF;
mem['h00FC] = 32'h03A00593;
mem['h00FD] = 32'h00C12503;
mem['h00FE] = 32'hCEDFF0EF;
mem['h00FF] = 32'h00812783;
mem['h0100] = 32'h00178793;
mem['h0101] = 32'h0007C783;
mem['h0102] = 32'h00200613;
mem['h0103] = 32'h00078593;
mem['h0104] = 32'h00C12503;
mem['h0105] = 32'hD39FF0EF;
mem['h0106] = 32'h03A00593;
mem['h0107] = 32'h00C12503;
mem['h0108] = 32'hCC5FF0EF;
mem['h0109] = 32'h00812783;
mem['h010A] = 32'h00278793;
mem['h010B] = 32'h0007C783;
mem['h010C] = 32'h00200613;
mem['h010D] = 32'h00078593;
mem['h010E] = 32'h00C12503;
mem['h010F] = 32'hD11FF0EF;
mem['h0110] = 32'h03A00593;
mem['h0111] = 32'h00C12503;
mem['h0112] = 32'hC9DFF0EF;
mem['h0113] = 32'h00812783;
mem['h0114] = 32'h00378793;
mem['h0115] = 32'h0007C783;
mem['h0116] = 32'h00200613;
mem['h0117] = 32'h00078593;
mem['h0118] = 32'h00C12503;
mem['h0119] = 32'hCE9FF0EF;
mem['h011A] = 32'h03A00593;
mem['h011B] = 32'h00C12503;
mem['h011C] = 32'hC75FF0EF;
mem['h011D] = 32'h00812783;
mem['h011E] = 32'h00478793;
mem['h011F] = 32'h0007C783;
mem['h0120] = 32'h00200613;
mem['h0121] = 32'h00078593;
mem['h0122] = 32'h00C12503;
mem['h0123] = 32'hCC1FF0EF;
mem['h0124] = 32'h03A00593;
mem['h0125] = 32'h00C12503;
mem['h0126] = 32'hC4DFF0EF;
mem['h0127] = 32'h00812783;
mem['h0128] = 32'h00578793;
mem['h0129] = 32'h0007C783;
mem['h012A] = 32'h00200613;
mem['h012B] = 32'h00078593;
mem['h012C] = 32'h00C12503;
mem['h012D] = 32'hC99FF0EF;
mem['h012E] = 32'h00000013;
mem['h012F] = 32'h01C12083;
mem['h0130] = 32'h02010113;
mem['h0131] = 32'h00008067;
mem['h0132] = 32'hFD010113;
mem['h0133] = 32'h02112623;
mem['h0134] = 32'h00A12623;
mem['h0135] = 32'h00B12423;
mem['h0136] = 32'h00C12783;
mem['h0137] = 32'h0047A783;
mem['h0138] = 32'h0007A783;
mem['h0139] = 32'h00078513;
mem['h013A] = 32'hB89FF0EF;
mem['h013B] = 32'h00A12E23;
mem['h013C] = 32'h01C12783;
mem['h013D] = 32'h1407D663;
mem['h013E] = 32'h01C12783;
mem['h013F] = 32'h0FF7F713;
mem['h0140] = 32'h01200793;
mem['h0141] = 32'h00F71663;
mem['h0142] = 32'h00000793;
mem['h0143] = 32'h1380006F;
mem['h0144] = 32'h00012C23;
mem['h0145] = 32'h1040006F;
mem['h0146] = 32'h01C12783;
mem['h0147] = 32'h0FF7F713;
mem['h0148] = 32'h00812783;
mem['h0149] = 32'h00E78023;
mem['h014A] = 32'h00812783;
mem['h014B] = 32'h0007C703;
mem['h014C] = 32'h00A00793;
mem['h014D] = 32'h0EF70A63;
mem['h014E] = 32'h00812783;
mem['h014F] = 32'h0007C703;
mem['h0150] = 32'h00D00793;
mem['h0151] = 32'h02F71063;
mem['h0152] = 32'h00D00593;
mem['h0153] = 32'h00C12503;
mem['h0154] = 32'hB95FF0EF;
mem['h0155] = 32'h00A00593;
mem['h0156] = 32'h00C12503;
mem['h0157] = 32'hB89FF0EF;
mem['h0158] = 32'h0CC0006F;
mem['h0159] = 32'h00812783;
mem['h015A] = 32'h0007C703;
mem['h015B] = 32'h00800793;
mem['h015C] = 32'h00F70A63;
mem['h015D] = 32'h00812783;
mem['h015E] = 32'h0007C703;
mem['h015F] = 32'h07F00793;
mem['h0160] = 32'h04F71663;
mem['h0161] = 32'h01812783;
mem['h0162] = 32'h06F05863;
mem['h0163] = 32'h00812783;
mem['h0164] = 32'hFFF78793;
mem['h0165] = 32'h00F12423;
mem['h0166] = 32'h01812783;
mem['h0167] = 32'hFFF78793;
mem['h0168] = 32'h00F12C23;
mem['h0169] = 32'h00800593;
mem['h016A] = 32'h00C12503;
mem['h016B] = 32'hB39FF0EF;
mem['h016C] = 32'h02000593;
mem['h016D] = 32'h00C12503;
mem['h016E] = 32'hB2DFF0EF;
mem['h016F] = 32'h00800593;
mem['h0170] = 32'h00C12503;
mem['h0171] = 32'hB21FF0EF;
mem['h0172] = 32'h0300006F;
mem['h0173] = 32'h00812783;
mem['h0174] = 32'h0007C783;
mem['h0175] = 32'h00078593;
mem['h0176] = 32'h00C12503;
mem['h0177] = 32'hB09FF0EF;
mem['h0178] = 32'h00812783;
mem['h0179] = 32'h00178793;
mem['h017A] = 32'h00F12423;
mem['h017B] = 32'h01812783;
mem['h017C] = 32'h00178793;
mem['h017D] = 32'h00F12C23;
mem['h017E] = 32'h00C12783;
mem['h017F] = 32'h0047A783;
mem['h0180] = 32'h0007A783;
mem['h0181] = 32'h00078513;
mem['h0182] = 32'hA69FF0EF;
mem['h0183] = 32'h00A12E23;
mem['h0184] = 32'h01C12783;
mem['h0185] = 32'hFE07D2E3;
mem['h0186] = 32'h01812703;
mem['h0187] = 32'h01E00793;
mem['h0188] = 32'hEEE7DCE3;
mem['h0189] = 32'h0080006F;
mem['h018A] = 32'h00000013;
mem['h018B] = 32'h00812783;
mem['h018C] = 32'h00078023;
mem['h018D] = 32'h01812783;
mem['h018E] = 32'h0FF7F793;
mem['h018F] = 32'h0080006F;
mem['h0190] = 32'h00000793;
mem['h0191] = 32'h00078513;
mem['h0192] = 32'h02C12083;
mem['h0193] = 32'h03010113;
mem['h0194] = 32'h00008067;
mem['h0195] = 32'hFB010113;
mem['h0196] = 32'h04112623;
mem['h0197] = 32'h00A12623;
mem['h0198] = 32'h000027B7;
mem['h0199] = 32'h65878793;
mem['h019A] = 32'h02F12C23;
mem['h019B] = 32'h000027B7;
mem['h019C] = 32'h66C78593;
mem['h019D] = 32'h00C12503;
mem['h019E] = 32'hC61FF0EF;
mem['h019F] = 32'h000027B7;
mem['h01A0] = 32'h68878593;
mem['h01A1] = 32'h00C12503;
mem['h01A2] = 32'hC51FF0EF;
mem['h01A3] = 32'h00300793;
mem['h01A4] = 32'h02F12E23;
mem['h01A5] = 32'h0D80006F;
mem['h01A6] = 32'h01410793;
mem['h01A7] = 32'h02F12A23;
mem['h01A8] = 32'h00000013;
mem['h01A9] = 32'h03412583;
mem['h01AA] = 32'h00C12503;
mem['h01AB] = 32'hE1DFF0EF;
mem['h01AC] = 32'h00050793;
mem['h01AD] = 32'h0017B793;
mem['h01AE] = 32'h0FF7F793;
mem['h01AF] = 32'hFE0794E3;
mem['h01B0] = 32'h000027B7;
mem['h01B1] = 32'h6C878593;
mem['h01B2] = 32'h00C12503;
mem['h01B3] = 32'hC0DFF0EF;
mem['h01B4] = 32'h03412583;
mem['h01B5] = 32'h00C12503;
mem['h01B6] = 32'hC01FF0EF;
mem['h01B7] = 32'h03412583;
mem['h01B8] = 32'h03812503;
mem['h01B9] = 32'h320010EF;
mem['h01BA] = 32'h00050793;
mem['h01BB] = 32'h0017B793;
mem['h01BC] = 32'h0FF7F793;
mem['h01BD] = 32'h00078C63;
mem['h01BE] = 32'h000027B7;
mem['h01BF] = 32'h6DC78593;
mem['h01C0] = 32'h00C12503;
mem['h01C1] = 32'hBD5FF0EF;
mem['h01C2] = 32'h06C0006F;
mem['h01C3] = 32'h000027B7;
mem['h01C4] = 32'h6F478593;
mem['h01C5] = 32'h00C12503;
mem['h01C6] = 32'hBC1FF0EF;
mem['h01C7] = 32'h03C12703;
mem['h01C8] = 32'h00100793;
mem['h01C9] = 32'h02E7DE63;
mem['h01CA] = 32'h000027B7;
mem['h01CB] = 32'h71078593;
mem['h01CC] = 32'h00C12503;
mem['h01CD] = 32'hBA5FF0EF;
mem['h01CE] = 32'h03C12783;
mem['h01CF] = 32'hFFF78793;
mem['h01D0] = 32'h00100613;
mem['h01D1] = 32'h00078593;
mem['h01D2] = 32'h00C12503;
mem['h01D3] = 32'hA01FF0EF;
mem['h01D4] = 32'h000027B7;
mem['h01D5] = 32'h73478593;
mem['h01D6] = 32'h00C12503;
mem['h01D7] = 32'hB7DFF0EF;
mem['h01D8] = 32'h03C12783;
mem['h01D9] = 32'hFFF78793;
mem['h01DA] = 32'h02F12E23;
mem['h01DB] = 32'h03C12783;
mem['h01DC] = 32'hF2F044E3;
mem['h01DD] = 32'h000027B7;
mem['h01DE] = 32'h73C78593;
mem['h01DF] = 32'h00C12503;
mem['h01E0] = 32'hB59FF0EF;
mem['h01E1] = 32'h00000013;
mem['h01E2] = 32'h04C12083;
mem['h01E3] = 32'h05010113;
mem['h01E4] = 32'h00008067;
mem['h01E5] = 32'hFF010113;
mem['h01E6] = 32'h00A12623;
mem['h01E7] = 32'h00B12423;
mem['h01E8] = 32'h00C12783;
mem['h01E9] = 32'h0007A783;
mem['h01EA] = 32'h0007A703;
mem['h01EB] = 32'h00077693;
mem['h01EC] = 32'h00812703;
mem['h01ED] = 32'h00E6E733;
mem['h01EE] = 32'h00E7A023;
mem['h01EF] = 32'h00000013;
mem['h01F0] = 32'h01010113;
mem['h01F1] = 32'h00008067;
mem['h01F2] = 32'hFF010113;
mem['h01F3] = 32'h00A12623;
mem['h01F4] = 32'h00B12423;
mem['h01F5] = 32'h00C12783;
mem['h01F6] = 32'h0007A783;
mem['h01F7] = 32'h0007A703;
mem['h01F8] = 32'h00077693;
mem['h01F9] = 32'h00812703;
mem['h01FA] = 32'h00E6E733;
mem['h01FB] = 32'h00E7A023;
mem['h01FC] = 32'h00000013;
mem['h01FD] = 32'h01010113;
mem['h01FE] = 32'h00008067;
mem['h01FF] = 32'hFF010113;
mem['h0200] = 32'h00A12623;
mem['h0201] = 32'h00B12423;
mem['h0202] = 32'h00C12783;
mem['h0203] = 32'h0007A783;
mem['h0204] = 32'h0007A703;
mem['h0205] = 32'h00077693;
mem['h0206] = 32'h00812703;
mem['h0207] = 32'h00E6E733;
mem['h0208] = 32'h00E7A023;
mem['h0209] = 32'h00000013;
mem['h020A] = 32'h01010113;
mem['h020B] = 32'h00008067;
mem['h020C] = 32'hFF010113;
mem['h020D] = 32'h00A12623;
mem['h020E] = 32'h00B12423;
mem['h020F] = 32'h00C12783;
mem['h0210] = 32'h0007A783;
mem['h0211] = 32'h0007A703;
mem['h0212] = 32'h00077693;
mem['h0213] = 32'h00812703;
mem['h0214] = 32'h00E6E733;
mem['h0215] = 32'h00E7A023;
mem['h0216] = 32'h00000013;
mem['h0217] = 32'h01010113;
mem['h0218] = 32'h00008067;
mem['h0219] = 32'hFF010113;
mem['h021A] = 32'h00A12623;
mem['h021B] = 32'h00B12423;
mem['h021C] = 32'h00C12783;
mem['h021D] = 32'h0007A783;
mem['h021E] = 32'h00812703;
mem['h021F] = 32'h00777713;
mem['h0220] = 32'h0FF77713;
mem['h0221] = 32'h00777713;
mem['h0222] = 32'h0007A683;
mem['h0223] = 32'hFF86F693;
mem['h0224] = 32'h00E6E733;
mem['h0225] = 32'h00E7A023;
mem['h0226] = 32'h00000013;
mem['h0227] = 32'h01010113;
mem['h0228] = 32'h00008067;
mem['h0229] = 32'hFF010113;
mem['h022A] = 32'h00A12623;
mem['h022B] = 32'h00B12423;
mem['h022C] = 32'h00C12783;
mem['h022D] = 32'h0007A783;
mem['h022E] = 32'h00812703;
mem['h022F] = 32'h00777713;
mem['h0230] = 32'h0FF77713;
mem['h0231] = 32'h00777713;
mem['h0232] = 32'h00371713;
mem['h0233] = 32'h0007A683;
mem['h0234] = 32'hFC76F693;
mem['h0235] = 32'h00E6E733;
mem['h0236] = 32'h00E7A023;
mem['h0237] = 32'h00000013;
mem['h0238] = 32'h01010113;
mem['h0239] = 32'h00008067;
mem['h023A] = 32'hFF010113;
mem['h023B] = 32'h00A12623;
mem['h023C] = 32'h00B12423;
mem['h023D] = 32'h00C12783;
mem['h023E] = 32'h0007A783;
mem['h023F] = 32'h00812703;
mem['h0240] = 32'h00177713;
mem['h0241] = 32'h0FF77713;
mem['h0242] = 32'h00177713;
mem['h0243] = 32'h00671713;
mem['h0244] = 32'h0007A683;
mem['h0245] = 32'hFBF6F693;
mem['h0246] = 32'h00E6E733;
mem['h0247] = 32'h00E7A023;
mem['h0248] = 32'h00000013;
mem['h0249] = 32'h01010113;
mem['h024A] = 32'h00008067;
mem['h024B] = 32'hFF010113;
mem['h024C] = 32'h00A12623;
mem['h024D] = 32'h00B12423;
mem['h024E] = 32'h00C12783;
mem['h024F] = 32'h0007A783;
mem['h0250] = 32'h00812703;
mem['h0251] = 32'h00177713;
mem['h0252] = 32'h0FF77713;
mem['h0253] = 32'h00177713;
mem['h0254] = 32'h00771713;
mem['h0255] = 32'h0007A683;
mem['h0256] = 32'hF7F6F693;
mem['h0257] = 32'h00E6E733;
mem['h0258] = 32'h00E7A023;
mem['h0259] = 32'h00000013;
mem['h025A] = 32'h01010113;
mem['h025B] = 32'h00008067;
mem['h025C] = 32'hFF010113;
mem['h025D] = 32'h00A12623;
mem['h025E] = 32'h00B12423;
mem['h025F] = 32'h00C12783;
mem['h0260] = 32'h0007A783;
mem['h0261] = 32'h00812703;
mem['h0262] = 32'h00177713;
mem['h0263] = 32'h0FF77713;
mem['h0264] = 32'h00177713;
mem['h0265] = 32'h00F71713;
mem['h0266] = 32'h0007A603;
mem['h0267] = 32'hFFFF86B7;
mem['h0268] = 32'hFFF68693;
mem['h0269] = 32'h00D676B3;
mem['h026A] = 32'h00E6E733;
mem['h026B] = 32'h00E7A023;
mem['h026C] = 32'h00000013;
mem['h026D] = 32'h01010113;
mem['h026E] = 32'h00008067;
mem['h026F] = 32'hFF010113;
mem['h0270] = 32'h00A12623;
mem['h0271] = 32'h00B12423;
mem['h0272] = 32'h00C12783;
mem['h0273] = 32'h0007A783;
mem['h0274] = 32'h00812703;
mem['h0275] = 32'h01071713;
mem['h0276] = 32'h01075713;
mem['h0277] = 32'h01071713;
mem['h0278] = 32'h0007A603;
mem['h0279] = 32'h000106B7;
mem['h027A] = 32'hFFF68693;
mem['h027B] = 32'h00D676B3;
mem['h027C] = 32'h00E6E733;
mem['h027D] = 32'h00E7A023;
mem['h027E] = 32'h00000013;
mem['h027F] = 32'h01010113;
mem['h0280] = 32'h00008067;
mem['h0281] = 32'hFF010113;
mem['h0282] = 32'h00A12623;
mem['h0283] = 32'h00B12423;
mem['h0284] = 32'h00C12783;
mem['h0285] = 32'h0007A783;
mem['h0286] = 32'h00812703;
mem['h0287] = 32'h00177713;
mem['h0288] = 32'h0FF77713;
mem['h0289] = 32'h00177713;
mem['h028A] = 32'h0007A683;
mem['h028B] = 32'hFFE6F693;
mem['h028C] = 32'h00E6E733;
mem['h028D] = 32'h00E7A023;
mem['h028E] = 32'h00000013;
mem['h028F] = 32'h01010113;
mem['h0290] = 32'h00008067;
mem['h0291] = 32'hFF010113;
mem['h0292] = 32'h00A12623;
mem['h0293] = 32'h00C12783;
mem['h0294] = 32'h0007A783;
mem['h0295] = 32'h0007A783;
mem['h0296] = 32'h0017F793;
mem['h0297] = 32'h0FF7F793;
mem['h0298] = 32'h00078513;
mem['h0299] = 32'h01010113;
mem['h029A] = 32'h00008067;
mem['h029B] = 32'hFF010113;
mem['h029C] = 32'h00A12623;
mem['h029D] = 32'h00C12783;
mem['h029E] = 32'h0007A783;
mem['h029F] = 32'h0007A783;
mem['h02A0] = 32'h00078513;
mem['h02A1] = 32'h01010113;
mem['h02A2] = 32'h00008067;
mem['h02A3] = 32'hFF010113;
mem['h02A4] = 32'h00A12623;
mem['h02A5] = 32'h00C12783;
mem['h02A6] = 32'h0007A783;
mem['h02A7] = 32'h0007A783;
mem['h02A8] = 32'h00078513;
mem['h02A9] = 32'h01010113;
mem['h02AA] = 32'h00008067;
mem['h02AB] = 32'hFF010113;
mem['h02AC] = 32'h00A12623;
mem['h02AD] = 32'h00C12783;
mem['h02AE] = 32'h0007A783;
mem['h02AF] = 32'h0007A783;
mem['h02B0] = 32'h00078513;
mem['h02B1] = 32'h01010113;
mem['h02B2] = 32'h00008067;
mem['h02B3] = 32'hFF010113;
mem['h02B4] = 32'h00A12623;
mem['h02B5] = 32'h00C12783;
mem['h02B6] = 32'h0007A783;
mem['h02B7] = 32'h0007A783;
mem['h02B8] = 32'h00078513;
mem['h02B9] = 32'h01010113;
mem['h02BA] = 32'h00008067;
mem['h02BB] = 32'hFF010113;
mem['h02BC] = 32'h00A12623;
mem['h02BD] = 32'h00C12783;
mem['h02BE] = 32'h0007A783;
mem['h02BF] = 32'h0007A783;
mem['h02C0] = 32'h0037D793;
mem['h02C1] = 32'h0077F793;
mem['h02C2] = 32'h0FF7F793;
mem['h02C3] = 32'h00078513;
mem['h02C4] = 32'h01010113;
mem['h02C5] = 32'h00008067;
mem['h02C6] = 32'hFF010113;
mem['h02C7] = 32'h00A12623;
mem['h02C8] = 32'h00C12783;
mem['h02C9] = 32'h0007A783;
mem['h02CA] = 32'h0007A783;
mem['h02CB] = 32'h00F7D793;
mem['h02CC] = 32'h0017F793;
mem['h02CD] = 32'h0FF7F793;
mem['h02CE] = 32'h00078513;
mem['h02CF] = 32'h01010113;
mem['h02D0] = 32'h00008067;
mem['h02D1] = 32'hFF010113;
mem['h02D2] = 32'h00A12623;
mem['h02D3] = 32'h00C12783;
mem['h02D4] = 32'h0007A783;
mem['h02D5] = 32'h0027D783;
mem['h02D6] = 32'h00078513;
mem['h02D7] = 32'h01010113;
mem['h02D8] = 32'h00008067;
mem['h02D9] = 32'hFF010113;
mem['h02DA] = 32'h00A12623;
mem['h02DB] = 32'h00B12423;
mem['h02DC] = 32'h00C12783;
mem['h02DD] = 32'h0007A783;
mem['h02DE] = 32'h00812703;
mem['h02DF] = 32'h00177713;
mem['h02E0] = 32'h0FF77713;
mem['h02E1] = 32'h00177713;
mem['h02E2] = 32'h0007A683;
mem['h02E3] = 32'hFFE6F693;
mem['h02E4] = 32'h00E6E733;
mem['h02E5] = 32'h00E7A023;
mem['h02E6] = 32'h00000013;
mem['h02E7] = 32'h01010113;
mem['h02E8] = 32'h00008067;
mem['h02E9] = 32'hFF010113;
mem['h02EA] = 32'h00A12623;
mem['h02EB] = 32'h00C12783;
mem['h02EC] = 32'h0007A783;
mem['h02ED] = 32'h0007A783;
mem['h02EE] = 32'h0017F793;
mem['h02EF] = 32'h0FF7F793;
mem['h02F0] = 32'h00078513;
mem['h02F1] = 32'h01010113;
mem['h02F2] = 32'h00008067;
mem['h02F3] = 32'hFD010113;
mem['h02F4] = 32'h02112623;
mem['h02F5] = 32'h00A12623;
mem['h02F6] = 32'h00B12423;
mem['h02F7] = 32'h00C12783;
mem['h02F8] = 32'h0007A783;
mem['h02F9] = 32'h0007A783;
mem['h02FA] = 32'h0187A783;
mem['h02FB] = 32'h00078513;
mem['h02FC] = 32'hE55FF0EF;
mem['h02FD] = 32'h00050793;
mem['h02FE] = 32'h00F037B3;
mem['h02FF] = 32'h0FF7F793;
mem['h0300] = 32'h26078063;
mem['h0301] = 32'h00012E23;
mem['h0302] = 32'h00C12783;
mem['h0303] = 32'h0007A783;
mem['h0304] = 32'h0007A783;
mem['h0305] = 32'h0107A703;
mem['h0306] = 32'h00812783;
mem['h0307] = 32'h0007C783;
mem['h0308] = 32'h00078593;
mem['h0309] = 32'h00070513;
mem['h030A] = 32'hC3DFF0EF;
mem['h030B] = 32'h00C12783;
mem['h030C] = 32'h0007A783;
mem['h030D] = 32'h0007A783;
mem['h030E] = 32'h0107A703;
mem['h030F] = 32'h00812783;
mem['h0310] = 32'h0017C783;
mem['h0311] = 32'h00078593;
mem['h0312] = 32'h00070513;
mem['h0313] = 32'hC59FF0EF;
mem['h0314] = 32'h00C12783;
mem['h0315] = 32'h0007A783;
mem['h0316] = 32'h0007A783;
mem['h0317] = 32'h0107A703;
mem['h0318] = 32'h00812783;
mem['h0319] = 32'h0027C783;
mem['h031A] = 32'h00078593;
mem['h031B] = 32'h00070513;
mem['h031C] = 32'hC79FF0EF;
mem['h031D] = 32'h00C12783;
mem['h031E] = 32'h0007A783;
mem['h031F] = 32'h0007A783;
mem['h0320] = 32'h0107A703;
mem['h0321] = 32'h00812783;
mem['h0322] = 32'h0037C783;
mem['h0323] = 32'h00078593;
mem['h0324] = 32'h00070513;
mem['h0325] = 32'hC99FF0EF;
mem['h0326] = 32'h00C12783;
mem['h0327] = 32'h0007A783;
mem['h0328] = 32'h0007A783;
mem['h0329] = 32'h0007A683;
mem['h032A] = 32'h00812783;
mem['h032B] = 32'h00878713;
mem['h032C] = 32'h01C12783;
mem['h032D] = 32'h00F707B3;
mem['h032E] = 32'h0007A783;
mem['h032F] = 32'h00078593;
mem['h0330] = 32'h00068513;
mem['h0331] = 32'hAD1FF0EF;
mem['h0332] = 32'h00C12783;
mem['h0333] = 32'h0007A783;
mem['h0334] = 32'h0007A783;
mem['h0335] = 32'h0047A683;
mem['h0336] = 32'h00812783;
mem['h0337] = 32'h00878713;
mem['h0338] = 32'h01C12783;
mem['h0339] = 32'h00478793;
mem['h033A] = 32'h00F707B3;
mem['h033B] = 32'h0007A783;
mem['h033C] = 32'h00078593;
mem['h033D] = 32'h00068513;
mem['h033E] = 32'hAD1FF0EF;
mem['h033F] = 32'h00C12783;
mem['h0340] = 32'h0007A783;
mem['h0341] = 32'h0007A783;
mem['h0342] = 32'h0087A683;
mem['h0343] = 32'h00812783;
mem['h0344] = 32'h00878713;
mem['h0345] = 32'h01C12783;
mem['h0346] = 32'h00878793;
mem['h0347] = 32'h00F707B3;
mem['h0348] = 32'h0007A783;
mem['h0349] = 32'h00078593;
mem['h034A] = 32'h00068513;
mem['h034B] = 32'hAD1FF0EF;
mem['h034C] = 32'h00C12783;
mem['h034D] = 32'h0007A783;
mem['h034E] = 32'h0007A783;
mem['h034F] = 32'h00C7A683;
mem['h0350] = 32'h00812783;
mem['h0351] = 32'h00878713;
mem['h0352] = 32'h01C12783;
mem['h0353] = 32'h00C78793;
mem['h0354] = 32'h00F707B3;
mem['h0355] = 32'h0007A783;
mem['h0356] = 32'h00078593;
mem['h0357] = 32'h00068513;
mem['h0358] = 32'hAD1FF0EF;
mem['h0359] = 32'h01C12783;
mem['h035A] = 32'h01078793;
mem['h035B] = 32'h00F12E23;
mem['h035C] = 32'h00812783;
mem['h035D] = 32'h0047A783;
mem['h035E] = 32'h01C12703;
mem['h035F] = 32'h06F77063;
mem['h0360] = 32'h00C12783;
mem['h0361] = 32'h0007A783;
mem['h0362] = 32'h0007A783;
mem['h0363] = 32'h0107A703;
mem['h0364] = 32'h000107B7;
mem['h0365] = 32'hFFF78593;
mem['h0366] = 32'h00070513;
mem['h0367] = 32'hC21FF0EF;
mem['h0368] = 32'h00C12783;
mem['h0369] = 32'h0007A783;
mem['h036A] = 32'h0007A783;
mem['h036B] = 32'h0107A783;
mem['h036C] = 32'h00000593;
mem['h036D] = 32'h00078513;
mem['h036E] = 32'hBB9FF0EF;
mem['h036F] = 32'h00C12783;
mem['h0370] = 32'h0007A783;
mem['h0371] = 32'h0007A783;
mem['h0372] = 32'h0147A783;
mem['h0373] = 32'h00100593;
mem['h0374] = 32'h00078513;
mem['h0375] = 32'hC31FF0EF;
mem['h0376] = 32'hEC1FF06F;
mem['h0377] = 32'h00812783;
mem['h0378] = 32'h0047A783;
mem['h0379] = 32'h01C12703;
mem['h037A] = 32'h40F707B3;
mem['h037B] = 32'h00F12C23;
mem['h037C] = 32'h00C12783;
mem['h037D] = 32'h0007A783;
mem['h037E] = 32'h0007A783;
mem['h037F] = 32'h0107A683;
mem['h0380] = 32'h01812783;
mem['h0381] = 32'h00010737;
mem['h0382] = 32'hFFF70713;
mem['h0383] = 32'h40F757B3;
mem['h0384] = 32'h00078593;
mem['h0385] = 32'h00068513;
mem['h0386] = 32'hBA5FF0EF;
mem['h0387] = 32'h00C12783;
mem['h0388] = 32'h0007A783;
mem['h0389] = 32'h0007A783;
mem['h038A] = 32'h0107A783;
mem['h038B] = 32'h00100593;
mem['h038C] = 32'h00078513;
mem['h038D] = 32'hB3DFF0EF;
mem['h038E] = 32'h00C12783;
mem['h038F] = 32'h0007A783;
mem['h0390] = 32'h0007A783;
mem['h0391] = 32'h0147A783;
mem['h0392] = 32'h00100593;
mem['h0393] = 32'h00078513;
mem['h0394] = 32'hBB5FF0EF;
mem['h0395] = 32'h00812783;
mem['h0396] = 32'h0047A783;
mem['h0397] = 32'h0080006F;
mem['h0398] = 32'h00000793;
mem['h0399] = 32'h00078513;
mem['h039A] = 32'h02C12083;
mem['h039B] = 32'h03010113;
mem['h039C] = 32'h00008067;
mem['h039D] = 32'hFD010113;
mem['h039E] = 32'h02112623;
mem['h039F] = 32'h02812423;
mem['h03A0] = 32'h00A12623;
mem['h03A1] = 32'h00B12423;
mem['h03A2] = 32'h00012E23;
mem['h03A3] = 32'h00812783;
mem['h03A4] = 32'h00078023;
mem['h03A5] = 32'h00812783;
mem['h03A6] = 32'h00078123;
mem['h03A7] = 32'h00812783;
mem['h03A8] = 32'h000781A3;
mem['h03A9] = 32'h00C12783;
mem['h03AA] = 32'h0007A783;
mem['h03AB] = 32'h0047A783;
mem['h03AC] = 32'h0187A783;
mem['h03AD] = 32'h00078513;
mem['h03AE] = 32'hCEDFF0EF;
mem['h03AF] = 32'h00050793;
mem['h03B0] = 32'h00F037B3;
mem['h03B1] = 32'h0FF7F793;
mem['h03B2] = 32'h1E078063;
mem['h03B3] = 32'h00C12783;
mem['h03B4] = 32'h0007A783;
mem['h03B5] = 32'h0047A783;
mem['h03B6] = 32'h0107A783;
mem['h03B7] = 32'h00078513;
mem['h03B8] = 32'hC0DFF0EF;
mem['h03B9] = 32'h00050793;
mem['h03BA] = 32'h0FF7F713;
mem['h03BB] = 32'h00812783;
mem['h03BC] = 32'h00E780A3;
mem['h03BD] = 32'h01C12703;
mem['h03BE] = 32'h5F000793;
mem['h03BF] = 32'h0CE7E863;
mem['h03C0] = 32'h00C12783;
mem['h03C1] = 32'h0007A783;
mem['h03C2] = 32'h0047A783;
mem['h03C3] = 32'h0007A683;
mem['h03C4] = 32'h00812783;
mem['h03C5] = 32'h00878713;
mem['h03C6] = 32'h01C12783;
mem['h03C7] = 32'h00F70433;
mem['h03C8] = 32'h00068513;
mem['h03C9] = 32'hB49FF0EF;
mem['h03CA] = 32'h00050793;
mem['h03CB] = 32'h00F42023;
mem['h03CC] = 32'h00C12783;
mem['h03CD] = 32'h0007A783;
mem['h03CE] = 32'h0047A783;
mem['h03CF] = 32'h0047A683;
mem['h03D0] = 32'h00812783;
mem['h03D1] = 32'h00878713;
mem['h03D2] = 32'h01C12783;
mem['h03D3] = 32'h00478793;
mem['h03D4] = 32'h00F70433;
mem['h03D5] = 32'h00068513;
mem['h03D6] = 32'hB35FF0EF;
mem['h03D7] = 32'h00050793;
mem['h03D8] = 32'h00F42023;
mem['h03D9] = 32'h00C12783;
mem['h03DA] = 32'h0007A783;
mem['h03DB] = 32'h0047A783;
mem['h03DC] = 32'h0087A683;
mem['h03DD] = 32'h00812783;
mem['h03DE] = 32'h00878713;
mem['h03DF] = 32'h01C12783;
mem['h03E0] = 32'h00878793;
mem['h03E1] = 32'h00F70433;
mem['h03E2] = 32'h00068513;
mem['h03E3] = 32'hB21FF0EF;
mem['h03E4] = 32'h00050793;
mem['h03E5] = 32'h00F42023;
mem['h03E6] = 32'h00C12783;
mem['h03E7] = 32'h0007A783;
mem['h03E8] = 32'h0047A783;
mem['h03E9] = 32'h00C7A683;
mem['h03EA] = 32'h00812783;
mem['h03EB] = 32'h00878713;
mem['h03EC] = 32'h01C12783;
mem['h03ED] = 32'h00C78793;
mem['h03EE] = 32'h00F70433;
mem['h03EF] = 32'h00068513;
mem['h03F0] = 32'hB0DFF0EF;
mem['h03F1] = 32'h00050793;
mem['h03F2] = 32'h00F42023;
mem['h03F3] = 32'h00C12783;
mem['h03F4] = 32'h0007A783;
mem['h03F5] = 32'h0047A783;
mem['h03F6] = 32'h0107A783;
mem['h03F7] = 32'h00078513;
mem['h03F8] = 32'hB39FF0EF;
mem['h03F9] = 32'h00050793;
mem['h03FA] = 32'h00F037B3;
mem['h03FB] = 32'h0FF7F793;
mem['h03FC] = 32'h08078663;
mem['h03FD] = 32'h00C12783;
mem['h03FE] = 32'h0007A783;
mem['h03FF] = 32'h0047A783;
mem['h0400] = 32'h0107A783;
mem['h0401] = 32'h00078513;
mem['h0402] = 32'hB3DFF0EF;
mem['h0403] = 32'h00050793;
mem['h0404] = 32'h00F11D23;
mem['h0405] = 32'h01C0006F;
mem['h0406] = 32'h01C12783;
mem['h0407] = 32'h00178793;
mem['h0408] = 32'h00F12E23;
mem['h0409] = 32'h01A15783;
mem['h040A] = 32'h0017D793;
mem['h040B] = 32'h00F11D23;
mem['h040C] = 32'h01A15783;
mem['h040D] = 32'h0017F793;
mem['h040E] = 32'hFE0790E3;
mem['h040F] = 32'h01C12783;
mem['h0410] = 32'h60000713;
mem['h0411] = 32'h00F77463;
mem['h0412] = 32'h60000793;
mem['h0413] = 32'h00812703;
mem['h0414] = 32'h00F72223;
mem['h0415] = 32'h00C12783;
mem['h0416] = 32'h0007A783;
mem['h0417] = 32'h0047A783;
mem['h0418] = 32'h0147A783;
mem['h0419] = 32'h00100593;
mem['h041A] = 32'h00078513;
mem['h041B] = 32'hAF9FF0EF;
mem['h041C] = 32'h00812783;
mem['h041D] = 32'h0047A783;
mem['h041E] = 32'h0340006F;
mem['h041F] = 32'h01C12783;
mem['h0420] = 32'h01078793;
mem['h0421] = 32'h00F12E23;
mem['h0422] = 32'h00C12783;
mem['h0423] = 32'h0007A783;
mem['h0424] = 32'h0047A783;
mem['h0425] = 32'h0147A783;
mem['h0426] = 32'h00100593;
mem['h0427] = 32'h00078513;
mem['h0428] = 32'hAC5FF0EF;
mem['h0429] = 32'hE51FF06F;
mem['h042A] = 32'h00000793;
mem['h042B] = 32'h00078513;
mem['h042C] = 32'h02C12083;
mem['h042D] = 32'h02812403;
mem['h042E] = 32'h03010113;
mem['h042F] = 32'h00008067;
mem['h0430] = 32'hFE010113;
mem['h0431] = 32'h00A12623;
mem['h0432] = 32'h00B12423;
mem['h0433] = 32'h00012E23;
mem['h0434] = 32'h00012C23;
mem['h0435] = 32'h0940006F;
mem['h0436] = 32'h00C12703;
mem['h0437] = 32'h01812783;
mem['h0438] = 32'h00F707B3;
mem['h0439] = 32'h0007C783;
mem['h043A] = 32'h01079793;
mem['h043B] = 32'h4107D793;
mem['h043C] = 32'h00879793;
mem['h043D] = 32'h01079713;
mem['h043E] = 32'h41075713;
mem['h043F] = 32'h01812783;
mem['h0440] = 32'h00178793;
mem['h0441] = 32'h00C12683;
mem['h0442] = 32'h00F687B3;
mem['h0443] = 32'h0007C783;
mem['h0444] = 32'h01079793;
mem['h0445] = 32'h4107D793;
mem['h0446] = 32'h00F767B3;
mem['h0447] = 32'h01079793;
mem['h0448] = 32'h4107D793;
mem['h0449] = 32'h00F11A23;
mem['h044A] = 32'h01415783;
mem['h044B] = 32'h01C12703;
mem['h044C] = 32'h00F707B3;
mem['h044D] = 32'h00F12E23;
mem['h044E] = 32'h01C12703;
mem['h044F] = 32'h000107B7;
mem['h0450] = 32'h00F76E63;
mem['h0451] = 32'h01C12703;
mem['h0452] = 32'h000107B7;
mem['h0453] = 32'hFFF78793;
mem['h0454] = 32'h00F777B3;
mem['h0455] = 32'h00178793;
mem['h0456] = 32'h00F12E23;
mem['h0457] = 32'h01812783;
mem['h0458] = 32'h00278793;
mem['h0459] = 32'h00F12C23;
mem['h045A] = 32'h01812783;
mem['h045B] = 32'h00178793;
mem['h045C] = 32'h00812703;
mem['h045D] = 32'hF6E7E2E3;
mem['h045E] = 32'h01812703;
mem['h045F] = 32'h00812783;
mem['h0460] = 32'h04F77863;
mem['h0461] = 32'h00C12703;
mem['h0462] = 32'h01812783;
mem['h0463] = 32'h00F707B3;
mem['h0464] = 32'h0007C783;
mem['h0465] = 32'h00879793;
mem['h0466] = 32'h00F11B23;
mem['h0467] = 32'h01615783;
mem['h0468] = 32'h01C12703;
mem['h0469] = 32'h00F707B3;
mem['h046A] = 32'h00F12E23;
mem['h046B] = 32'h01C12703;
mem['h046C] = 32'h000107B7;
mem['h046D] = 32'h00F76E63;
mem['h046E] = 32'h01C12703;
mem['h046F] = 32'h000107B7;
mem['h0470] = 32'hFFF78793;
mem['h0471] = 32'h00F777B3;
mem['h0472] = 32'h00178793;
mem['h0473] = 32'h00F12E23;
mem['h0474] = 32'h01C12783;
mem['h0475] = 32'h01079793;
mem['h0476] = 32'h0107D793;
mem['h0477] = 32'hFFF7C793;
mem['h0478] = 32'h01079793;
mem['h0479] = 32'h0107D793;
mem['h047A] = 32'h00078513;
mem['h047B] = 32'h02010113;
mem['h047C] = 32'h00008067;
mem['h047D] = 32'hFE010113;
mem['h047E] = 32'h00A12623;
mem['h047F] = 32'h00C12783;
mem['h0480] = 32'h00878793;
mem['h0481] = 32'h00F12E23;
mem['h0482] = 32'h00C12783;
mem['h0483] = 32'h00878793;
mem['h0484] = 32'h00E78793;
mem['h0485] = 32'h00F12C23;
mem['h0486] = 32'h01C12783;
mem['h0487] = 32'h00C7C703;
mem['h0488] = 32'h00800793;
mem['h0489] = 32'h00F71E63;
mem['h048A] = 32'h01C12783;
mem['h048B] = 32'h00D7C703;
mem['h048C] = 32'h00600793;
mem['h048D] = 32'h00F71663;
mem['h048E] = 32'h00100793;
mem['h048F] = 32'h06C0006F;
mem['h0490] = 32'h01C12783;
mem['h0491] = 32'h00C7C703;
mem['h0492] = 32'h00800793;
mem['h0493] = 32'h04F71C63;
mem['h0494] = 32'h01C12783;
mem['h0495] = 32'h00D7C783;
mem['h0496] = 32'h04079663;
mem['h0497] = 32'h01812783;
mem['h0498] = 32'h0007C783;
mem['h0499] = 32'hFF07F793;
mem['h049A] = 32'h0FF7F713;
mem['h049B] = 32'h04000793;
mem['h049C] = 32'h02F71A63;
mem['h049D] = 32'h01812783;
mem['h049E] = 32'h0097C703;
mem['h049F] = 32'h00100793;
mem['h04A0] = 32'h00F71663;
mem['h04A1] = 32'h00200793;
mem['h04A2] = 32'h0200006F;
mem['h04A3] = 32'h01812783;
mem['h04A4] = 32'h0097C703;
mem['h04A5] = 32'h01100793;
mem['h04A6] = 32'h00F71663;
mem['h04A7] = 32'h00300793;
mem['h04A8] = 32'h0080006F;
mem['h04A9] = 32'h00000793;
mem['h04AA] = 32'h00078513;
mem['h04AB] = 32'h02010113;
mem['h04AC] = 32'h00008067;
mem['h04AD] = 32'hFD010113;
mem['h04AE] = 32'h02112623;
mem['h04AF] = 32'h00A12623;
mem['h04B0] = 32'h00B12423;
mem['h04B1] = 32'h00C12223;
mem['h04B2] = 32'h00D12023;
mem['h04B3] = 32'h00412783;
mem['h04B4] = 32'h00878793;
mem['h04B5] = 32'h00F12E23;
mem['h04B6] = 32'h00412783;
mem['h04B7] = 32'h00878793;
mem['h04B8] = 32'h00E78793;
mem['h04B9] = 32'h00F12C23;
mem['h04BA] = 32'h00012783;
mem['h04BB] = 32'h00878793;
mem['h04BC] = 32'h00F12A23;
mem['h04BD] = 32'h00012783;
mem['h04BE] = 32'h00878793;
mem['h04BF] = 32'h00E78793;
mem['h04C0] = 32'h00F12823;
mem['h04C1] = 32'h01812783;
mem['h04C2] = 32'h0007C783;
mem['h04C3] = 32'h00079A63;
mem['h04C4] = 32'h01812783;
mem['h04C5] = 32'h0017C703;
mem['h04C6] = 32'h00100793;
mem['h04C7] = 32'h00F70663;
mem['h04C8] = 32'h00000793;
mem['h04C9] = 32'h1D00006F;
mem['h04CA] = 32'h01812783;
mem['h04CB] = 32'h0027C703;
mem['h04CC] = 32'h00800793;
mem['h04CD] = 32'h00F71863;
mem['h04CE] = 32'h01812783;
mem['h04CF] = 32'h0037C783;
mem['h04D0] = 32'h00078663;
mem['h04D1] = 32'h00000793;
mem['h04D2] = 32'h1AC0006F;
mem['h04D3] = 32'h01812783;
mem['h04D4] = 32'h01878793;
mem['h04D5] = 32'h00C12703;
mem['h04D6] = 32'h00400613;
mem['h04D7] = 32'h00070593;
mem['h04D8] = 32'h00078513;
mem['h04D9] = 32'h5C0000EF;
mem['h04DA] = 32'h00050793;
mem['h04DB] = 32'h00F037B3;
mem['h04DC] = 32'h0FF7F793;
mem['h04DD] = 32'h00078663;
mem['h04DE] = 32'h00000793;
mem['h04DF] = 32'h1780006F;
mem['h04E0] = 32'h01812783;
mem['h04E1] = 32'h0067C783;
mem['h04E2] = 32'h16079463;
mem['h04E3] = 32'h01812783;
mem['h04E4] = 32'h0077C703;
mem['h04E5] = 32'h00100793;
mem['h04E6] = 32'h14F71C63;
mem['h04E7] = 32'h00412783;
mem['h04E8] = 32'h0017C703;
mem['h04E9] = 32'h00012783;
mem['h04EA] = 32'h00E78023;
mem['h04EB] = 32'h00012783;
mem['h04EC] = 32'h00100713;
mem['h04ED] = 32'h00E781A3;
mem['h04EE] = 32'h00012783;
mem['h04EF] = 32'h02A00713;
mem['h04F0] = 32'h00E7A223;
mem['h04F1] = 32'h01412703;
mem['h04F2] = 32'h01812783;
mem['h04F3] = 32'h00878793;
mem['h04F4] = 32'h00600613;
mem['h04F5] = 32'h00078593;
mem['h04F6] = 32'h00070513;
mem['h04F7] = 32'h4D8000EF;
mem['h04F8] = 32'h01412783;
mem['h04F9] = 32'h00678713;
mem['h04FA] = 32'h00C12783;
mem['h04FB] = 32'h00878793;
mem['h04FC] = 32'h00600613;
mem['h04FD] = 32'h00078593;
mem['h04FE] = 32'h00070513;
mem['h04FF] = 32'h4B8000EF;
mem['h0500] = 32'h01412783;
mem['h0501] = 32'h00800713;
mem['h0502] = 32'h00E78623;
mem['h0503] = 32'h01412783;
mem['h0504] = 32'h00600713;
mem['h0505] = 32'h00E786A3;
mem['h0506] = 32'h01012783;
mem['h0507] = 32'h00078023;
mem['h0508] = 32'h01012783;
mem['h0509] = 32'h00100713;
mem['h050A] = 32'h00E780A3;
mem['h050B] = 32'h01012783;
mem['h050C] = 32'h00800713;
mem['h050D] = 32'h00E78123;
mem['h050E] = 32'h01012783;
mem['h050F] = 32'h000781A3;
mem['h0510] = 32'h01012783;
mem['h0511] = 32'h00600713;
mem['h0512] = 32'h00E78223;
mem['h0513] = 32'h01012783;
mem['h0514] = 32'h00400713;
mem['h0515] = 32'h00E782A3;
mem['h0516] = 32'h01012783;
mem['h0517] = 32'h00078323;
mem['h0518] = 32'h01012783;
mem['h0519] = 32'h00200713;
mem['h051A] = 32'h00E783A3;
mem['h051B] = 32'h01012783;
mem['h051C] = 32'h00878713;
mem['h051D] = 32'h00C12783;
mem['h051E] = 32'h00878793;
mem['h051F] = 32'h00600613;
mem['h0520] = 32'h00078593;
mem['h0521] = 32'h00070513;
mem['h0522] = 32'h42C000EF;
mem['h0523] = 32'h01012783;
mem['h0524] = 32'h00E78793;
mem['h0525] = 32'h00C12703;
mem['h0526] = 32'h00400613;
mem['h0527] = 32'h00070593;
mem['h0528] = 32'h00078513;
mem['h0529] = 32'h410000EF;
mem['h052A] = 32'h01012783;
mem['h052B] = 32'h01278713;
mem['h052C] = 32'h01812783;
mem['h052D] = 32'h00878793;
mem['h052E] = 32'h00600613;
mem['h052F] = 32'h00078593;
mem['h0530] = 32'h00070513;
mem['h0531] = 32'h3F0000EF;
mem['h0532] = 32'h01012783;
mem['h0533] = 32'h01878713;
mem['h0534] = 32'h01812783;
mem['h0535] = 32'h00E78793;
mem['h0536] = 32'h00400613;
mem['h0537] = 32'h00078593;
mem['h0538] = 32'h00070513;
mem['h0539] = 32'h3D0000EF;
mem['h053A] = 32'h00100793;
mem['h053B] = 32'h0080006F;
mem['h053C] = 32'h00000793;
mem['h053D] = 32'h00078513;
mem['h053E] = 32'h02C12083;
mem['h053F] = 32'h03010113;
mem['h0540] = 32'h00008067;
mem['h0541] = 32'hFC010113;
mem['h0542] = 32'h02112E23;
mem['h0543] = 32'h00A12623;
mem['h0544] = 32'h00B12423;
mem['h0545] = 32'h00C12223;
mem['h0546] = 32'h00812783;
mem['h0547] = 32'h00878793;
mem['h0548] = 32'h02F12623;
mem['h0549] = 32'h00812783;
mem['h054A] = 32'h00878793;
mem['h054B] = 32'h00E78793;
mem['h054C] = 32'h02F12423;
mem['h054D] = 32'h00812783;
mem['h054E] = 32'h00878793;
mem['h054F] = 32'h02278793;
mem['h0550] = 32'h02F12223;
mem['h0551] = 32'h00412783;
mem['h0552] = 32'h00878793;
mem['h0553] = 32'h02F12023;
mem['h0554] = 32'h00412783;
mem['h0555] = 32'h00878793;
mem['h0556] = 32'h00E78793;
mem['h0557] = 32'h00F12E23;
mem['h0558] = 32'h00412783;
mem['h0559] = 32'h00878793;
mem['h055A] = 32'h02278793;
mem['h055B] = 32'h00F12C23;
mem['h055C] = 32'h02812783;
mem['h055D] = 32'h01078793;
mem['h055E] = 32'h00C12703;
mem['h055F] = 32'h00400613;
mem['h0560] = 32'h00070593;
mem['h0561] = 32'h00078513;
mem['h0562] = 32'h39C000EF;
mem['h0563] = 32'h00050793;
mem['h0564] = 32'h00F037B3;
mem['h0565] = 32'h0FF7F793;
mem['h0566] = 32'h00078663;
mem['h0567] = 32'h00000793;
mem['h0568] = 32'h2A00006F;
mem['h0569] = 32'h02412783;
mem['h056A] = 32'h0007C703;
mem['h056B] = 32'h00800793;
mem['h056C] = 32'h28F71663;
mem['h056D] = 32'h02412783;
mem['h056E] = 32'h0017C783;
mem['h056F] = 32'h28079063;
mem['h0570] = 32'h00812783;
mem['h0571] = 32'h0017C703;
mem['h0572] = 32'h00412783;
mem['h0573] = 32'h00E78023;
mem['h0574] = 32'h00412783;
mem['h0575] = 32'h00100713;
mem['h0576] = 32'h00E781A3;
mem['h0577] = 32'h00812783;
mem['h0578] = 32'h0047A703;
mem['h0579] = 32'h00412783;
mem['h057A] = 32'h00E7A223;
mem['h057B] = 32'h02012703;
mem['h057C] = 32'h02C12783;
mem['h057D] = 32'h00678793;
mem['h057E] = 32'h00600613;
mem['h057F] = 32'h00078593;
mem['h0580] = 32'h00070513;
mem['h0581] = 32'h2B0000EF;
mem['h0582] = 32'h02012783;
mem['h0583] = 32'h00678713;
mem['h0584] = 32'h00C12783;
mem['h0585] = 32'h00878793;
mem['h0586] = 32'h00600613;
mem['h0587] = 32'h00078593;
mem['h0588] = 32'h00070513;
mem['h0589] = 32'h290000EF;
mem['h058A] = 32'h02012783;
mem['h058B] = 32'h00800713;
mem['h058C] = 32'h00E78623;
mem['h058D] = 32'h02012783;
mem['h058E] = 32'h000786A3;
mem['h058F] = 32'h01C12783;
mem['h0590] = 32'h0007C703;
mem['h0591] = 32'hFF077713;
mem['h0592] = 32'h00576713;
mem['h0593] = 32'h00E78023;
mem['h0594] = 32'h01C12783;
mem['h0595] = 32'h0007C703;
mem['h0596] = 32'h00F77713;
mem['h0597] = 32'h04076713;
mem['h0598] = 32'h00E78023;
mem['h0599] = 32'h01C12783;
mem['h059A] = 32'h000780A3;
mem['h059B] = 32'h02812783;
mem['h059C] = 32'h0027C703;
mem['h059D] = 32'h01C12783;
mem['h059E] = 32'h00E78123;
mem['h059F] = 32'h02812783;
mem['h05A0] = 32'h0037C703;
mem['h05A1] = 32'h01C12783;
mem['h05A2] = 32'h00E781A3;
mem['h05A3] = 32'h01C12783;
mem['h05A4] = 32'h00078223;
mem['h05A5] = 32'h01C12783;
mem['h05A6] = 32'h000782A3;
mem['h05A7] = 32'h01C12783;
mem['h05A8] = 32'h00079323;
mem['h05A9] = 32'h01C12783;
mem['h05AA] = 32'hFFF00713;
mem['h05AB] = 32'h00E78423;
mem['h05AC] = 32'h01C12783;
mem['h05AD] = 32'h00100713;
mem['h05AE] = 32'h00E784A3;
mem['h05AF] = 32'h01C12783;
mem['h05B0] = 32'h00078523;
mem['h05B1] = 32'h01C12783;
mem['h05B2] = 32'h000785A3;
mem['h05B3] = 32'h01C12783;
mem['h05B4] = 32'h00C78793;
mem['h05B5] = 32'h00C12703;
mem['h05B6] = 32'h00400613;
mem['h05B7] = 32'h00070593;
mem['h05B8] = 32'h00078513;
mem['h05B9] = 32'h1D0000EF;
mem['h05BA] = 32'h01C12783;
mem['h05BB] = 32'h01078713;
mem['h05BC] = 32'h02812783;
mem['h05BD] = 32'h00C78793;
mem['h05BE] = 32'h00400613;
mem['h05BF] = 32'h00078593;
mem['h05C0] = 32'h00070513;
mem['h05C1] = 32'h1B0000EF;
mem['h05C2] = 32'h00412783;
mem['h05C3] = 32'h00878793;
mem['h05C4] = 32'h00E78793;
mem['h05C5] = 32'h01400593;
mem['h05C6] = 32'h00078513;
mem['h05C7] = 32'h9A5FF0EF;
mem['h05C8] = 32'h00050793;
mem['h05C9] = 32'h00F11B23;
mem['h05CA] = 32'h01615783;
mem['h05CB] = 32'h0087D793;
mem['h05CC] = 32'h01079793;
mem['h05CD] = 32'h0107D793;
mem['h05CE] = 32'h0FF7F713;
mem['h05CF] = 32'h01C12783;
mem['h05D0] = 32'h00E78523;
mem['h05D1] = 32'h01615783;
mem['h05D2] = 32'h0FF7F713;
mem['h05D3] = 32'h01C12783;
mem['h05D4] = 32'h00E785A3;
mem['h05D5] = 32'h01812783;
mem['h05D6] = 32'h00078023;
mem['h05D7] = 32'h01812783;
mem['h05D8] = 32'h000780A3;
mem['h05D9] = 32'h01812783;
mem['h05DA] = 32'h00078123;
mem['h05DB] = 32'h01812783;
mem['h05DC] = 32'h000781A3;
mem['h05DD] = 32'h02412783;
mem['h05DE] = 32'h0047C703;
mem['h05DF] = 32'h01812783;
mem['h05E0] = 32'h00E78223;
mem['h05E1] = 32'h02412783;
mem['h05E2] = 32'h0057C703;
mem['h05E3] = 32'h01812783;
mem['h05E4] = 32'h00E782A3;
mem['h05E5] = 32'h02412783;
mem['h05E6] = 32'h0067C703;
mem['h05E7] = 32'h01812783;
mem['h05E8] = 32'h00E78323;
mem['h05E9] = 32'h02412783;
mem['h05EA] = 32'h0077C703;
mem['h05EB] = 32'h01812783;
mem['h05EC] = 32'h00E783A3;
mem['h05ED] = 32'h00412783;
mem['h05EE] = 32'h00878793;
mem['h05EF] = 32'h02A78713;
mem['h05F0] = 32'h00812783;
mem['h05F1] = 32'h00878793;
mem['h05F2] = 32'h02A78693;
mem['h05F3] = 32'h00812783;
mem['h05F4] = 32'h0047A783;
mem['h05F5] = 32'hFD678793;
mem['h05F6] = 32'h00078613;
mem['h05F7] = 32'h00068593;
mem['h05F8] = 32'h00070513;
mem['h05F9] = 32'h0D0000EF;
mem['h05FA] = 32'h00812783;
mem['h05FB] = 32'h0047A783;
mem['h05FC] = 32'hFDE78793;
mem['h05FD] = 32'h00078593;
mem['h05FE] = 32'h01812503;
mem['h05FF] = 32'h8C5FF0EF;
mem['h0600] = 32'h00050793;
mem['h0601] = 32'h00F11B23;
mem['h0602] = 32'h01615783;
mem['h0603] = 32'h0087D793;
mem['h0604] = 32'h01079793;
mem['h0605] = 32'h0107D793;
mem['h0606] = 32'h0FF7F713;
mem['h0607] = 32'h01812783;
mem['h0608] = 32'h00E78123;
mem['h0609] = 32'h01615783;
mem['h060A] = 32'h0FF7F713;
mem['h060B] = 32'h01812783;
mem['h060C] = 32'h00E781A3;
mem['h060D] = 32'h00100793;
mem['h060E] = 32'h0080006F;
mem['h060F] = 32'h00000793;
mem['h0610] = 32'h00078513;
mem['h0611] = 32'h03C12083;
mem['h0612] = 32'h04010113;
mem['h0613] = 32'h00008067;
mem['h0614] = 32'hFE010113;
mem['h0615] = 32'h00A12623;
mem['h0616] = 32'h00B12423;
mem['h0617] = 32'h00C12223;
mem['h0618] = 32'h00C12783;
mem['h0619] = 32'h00F12C23;
mem['h061A] = 32'h00812783;
mem['h061B] = 32'h00F10BA3;
mem['h061C] = 32'h00012E23;
mem['h061D] = 32'h0240006F;
mem['h061E] = 32'h01812703;
mem['h061F] = 32'h01C12783;
mem['h0620] = 32'h00F707B3;
mem['h0621] = 32'h01714703;
mem['h0622] = 32'h00E78023;
mem['h0623] = 32'h01C12783;
mem['h0624] = 32'h00178793;
mem['h0625] = 32'h00F12E23;
mem['h0626] = 32'h01C12703;
mem['h0627] = 32'h00412783;
mem['h0628] = 32'hFCF76CE3;
mem['h0629] = 32'h00C12783;
mem['h062A] = 32'h00078513;
mem['h062B] = 32'h02010113;
mem['h062C] = 32'h00008067;
mem['h062D] = 32'hFE010113;
mem['h062E] = 32'h00A12623;
mem['h062F] = 32'h00B12423;
mem['h0630] = 32'h00C12223;
mem['h0631] = 32'h00C12783;
mem['h0632] = 32'h00F12C23;
mem['h0633] = 32'h00812783;
mem['h0634] = 32'h00F12A23;
mem['h0635] = 32'h00012E23;
mem['h0636] = 32'h0300006F;
mem['h0637] = 32'h01412703;
mem['h0638] = 32'h01C12783;
mem['h0639] = 32'h00F70733;
mem['h063A] = 32'h01812683;
mem['h063B] = 32'h01C12783;
mem['h063C] = 32'h00F687B3;
mem['h063D] = 32'h00074703;
mem['h063E] = 32'h00E78023;
mem['h063F] = 32'h01C12783;
mem['h0640] = 32'h00178793;
mem['h0641] = 32'h00F12E23;
mem['h0642] = 32'h01C12703;
mem['h0643] = 32'h00412783;
mem['h0644] = 32'hFCF766E3;
mem['h0645] = 32'h00C12783;
mem['h0646] = 32'h00078513;
mem['h0647] = 32'h02010113;
mem['h0648] = 32'h00008067;
mem['h0649] = 32'hFE010113;
mem['h064A] = 32'h00A12623;
mem['h064B] = 32'h00B12423;
mem['h064C] = 32'h00C12223;
mem['h064D] = 32'h00C12783;
mem['h064E] = 32'h00F12C23;
mem['h064F] = 32'h00812783;
mem['h0650] = 32'h00F12A23;
mem['h0651] = 32'h00012E23;
mem['h0652] = 32'h0600006F;
mem['h0653] = 32'h01812703;
mem['h0654] = 32'h01C12783;
mem['h0655] = 32'h00F707B3;
mem['h0656] = 32'h0007C703;
mem['h0657] = 32'h01412683;
mem['h0658] = 32'h01C12783;
mem['h0659] = 32'h00F687B3;
mem['h065A] = 32'h0007C783;
mem['h065B] = 32'h02F70863;
mem['h065C] = 32'h01812703;
mem['h065D] = 32'h01C12783;
mem['h065E] = 32'h00F707B3;
mem['h065F] = 32'h0007C783;
mem['h0660] = 32'h00078693;
mem['h0661] = 32'h01412703;
mem['h0662] = 32'h01C12783;
mem['h0663] = 32'h00F707B3;
mem['h0664] = 32'h0007C783;
mem['h0665] = 32'h40F687B3;
mem['h0666] = 32'h0200006F;
mem['h0667] = 32'h01C12783;
mem['h0668] = 32'h00178793;
mem['h0669] = 32'h00F12E23;
mem['h066A] = 32'h01C12703;
mem['h066B] = 32'h00412783;
mem['h066C] = 32'hF8F76EE3;
mem['h066D] = 32'h00000793;
mem['h066E] = 32'h00078513;
mem['h066F] = 32'h02010113;
mem['h0670] = 32'h00008067;
mem['h0671] = 32'hFE010113;
mem['h0672] = 32'h00A12623;
mem['h0673] = 32'h00012E23;
mem['h0674] = 32'h0100006F;
mem['h0675] = 32'h01C12783;
mem['h0676] = 32'h00178793;
mem['h0677] = 32'h00F12E23;
mem['h0678] = 32'h00C12703;
mem['h0679] = 32'h01C12783;
mem['h067A] = 32'h00F707B3;
mem['h067B] = 32'h0007C783;
mem['h067C] = 32'hFE0792E3;
mem['h067D] = 32'h01C12783;
mem['h067E] = 32'h00078513;
mem['h067F] = 32'h02010113;
mem['h0680] = 32'h00008067;
mem['h0681] = 32'hFE010113;
mem['h0682] = 32'h00112E23;
mem['h0683] = 32'h00A12623;
mem['h0684] = 32'h00B12423;
mem['h0685] = 32'h00C12503;
mem['h0686] = 32'hFADFF0EF;
mem['h0687] = 32'h00050793;
mem['h0688] = 32'h00078613;
mem['h0689] = 32'h00812583;
mem['h068A] = 32'h00C12503;
mem['h068B] = 32'hEF9FF0EF;
mem['h068C] = 32'h00050793;
mem['h068D] = 32'h00078513;
mem['h068E] = 32'h01C12083;
mem['h068F] = 32'h02010113;
mem['h0690] = 32'h00008067;
mem['h0691] = 32'hFE010113;
mem['h0692] = 32'h00A12623;
mem['h0693] = 32'h0001A783;
mem['h0694] = 32'h00078713;
mem['h0695] = 32'h100007B7;
mem['h0696] = 32'h00078793;
mem['h0697] = 32'h00F707B3;
mem['h0698] = 32'h00F12E23;
mem['h0699] = 32'h0001A703;
mem['h069A] = 32'h00C12783;
mem['h069B] = 32'h00F70733;
mem['h069C] = 32'h00E1A023;
mem['h069D] = 32'h0001A703;
mem['h069E] = 32'h000017B7;
mem['h069F] = 32'h80078793;
mem['h06A0] = 32'h00E7D463;
mem['h06A1] = 32'h00100073;
mem['h06A2] = 32'h01C12783;
mem['h06A3] = 32'h00078513;
mem['h06A4] = 32'h02010113;
mem['h06A5] = 32'h00008067;
mem['h06A6] = 32'hFE010113;
mem['h06A7] = 32'h00112E23;
mem['h06A8] = 32'h00A12623;
mem['h06A9] = 32'h00C12783;
mem['h06AA] = 32'h00078513;
mem['h06AB] = 32'hF99FF0EF;
mem['h06AC] = 32'h00050793;
mem['h06AD] = 32'h00078513;
mem['h06AE] = 32'h01C12083;
mem['h06AF] = 32'h02010113;
mem['h06B0] = 32'h00008067;
mem['h06B1] = 32'hFF010113;
mem['h06B2] = 32'h00A12623;
mem['h06B3] = 32'h00000013;
mem['h06B4] = 32'h01010113;
mem['h06B5] = 32'h00008067;
mem['h06B6] = 32'hFF010113;
mem['h06B7] = 32'h00A12623;
mem['h06B8] = 32'h00B12423;
mem['h06B9] = 32'h00C12783;
mem['h06BA] = 32'h00812703;
mem['h06BB] = 32'h00E7A023;
mem['h06BC] = 32'h00000013;
mem['h06BD] = 32'h01010113;
mem['h06BE] = 32'h00008067;
mem['h06BF] = 32'hFF010113;
mem['h06C0] = 32'h00A12623;
mem['h06C1] = 32'h00B12423;
mem['h06C2] = 32'h00C12783;
mem['h06C3] = 32'h00812703;
mem['h06C4] = 32'h00E7A023;
mem['h06C5] = 32'h00000013;
mem['h06C6] = 32'h01010113;
mem['h06C7] = 32'h00008067;
mem['h06C8] = 32'hFF010113;
mem['h06C9] = 32'h00A12623;
mem['h06CA] = 32'h00B12423;
mem['h06CB] = 32'h00C12783;
mem['h06CC] = 32'h00812703;
mem['h06CD] = 32'h00E7A023;
mem['h06CE] = 32'h00000013;
mem['h06CF] = 32'h01010113;
mem['h06D0] = 32'h00008067;
mem['h06D1] = 32'hFF010113;
mem['h06D2] = 32'h00A12623;
mem['h06D3] = 32'h00B12423;
mem['h06D4] = 32'h00C12783;
mem['h06D5] = 32'h00812703;
mem['h06D6] = 32'h00E7A023;
mem['h06D7] = 32'h00000013;
mem['h06D8] = 32'h01010113;
mem['h06D9] = 32'h00008067;
mem['h06DA] = 32'hFF010113;
mem['h06DB] = 32'h00A12623;
mem['h06DC] = 32'h00B12423;
mem['h06DD] = 32'h00C12783;
mem['h06DE] = 32'h00812703;
mem['h06DF] = 32'h00E7A023;
mem['h06E0] = 32'h00000013;
mem['h06E1] = 32'h01010113;
mem['h06E2] = 32'h00008067;
mem['h06E3] = 32'hFF010113;
mem['h06E4] = 32'h00A12623;
mem['h06E5] = 32'h00B12423;
mem['h06E6] = 32'h00C12783;
mem['h06E7] = 32'h00812703;
mem['h06E8] = 32'h00E7A023;
mem['h06E9] = 32'h00000013;
mem['h06EA] = 32'h01010113;
mem['h06EB] = 32'h00008067;
mem['h06EC] = 32'hFF010113;
mem['h06ED] = 32'h00A12623;
mem['h06EE] = 32'h00B12423;
mem['h06EF] = 32'h00C12783;
mem['h06F0] = 32'h00812703;
mem['h06F1] = 32'h00E7A023;
mem['h06F2] = 32'h00000013;
mem['h06F3] = 32'h01010113;
mem['h06F4] = 32'h00008067;
mem['h06F5] = 32'hFE010113;
mem['h06F6] = 32'h00112E23;
mem['h06F7] = 32'h00812C23;
mem['h06F8] = 32'h00A12623;
mem['h06F9] = 32'h00B12423;
mem['h06FA] = 32'h00400513;
mem['h06FB] = 32'hEADFF0EF;
mem['h06FC] = 32'h00050793;
mem['h06FD] = 32'h00078413;
mem['h06FE] = 32'h00812583;
mem['h06FF] = 32'h00040513;
mem['h0700] = 32'hED9FF0EF;
mem['h0701] = 32'h00C12783;
mem['h0702] = 32'h0087A023;
mem['h0703] = 32'h00400513;
mem['h0704] = 32'hE89FF0EF;
mem['h0705] = 32'h00050793;
mem['h0706] = 32'h00078413;
mem['h0707] = 32'h00812783;
mem['h0708] = 32'h00478793;
mem['h0709] = 32'h00078593;
mem['h070A] = 32'h00040513;
mem['h070B] = 32'hED1FF0EF;
mem['h070C] = 32'h00C12783;
mem['h070D] = 32'h0087A223;
mem['h070E] = 32'h00400513;
mem['h070F] = 32'hE5DFF0EF;
mem['h0710] = 32'h00050793;
mem['h0711] = 32'h00078413;
mem['h0712] = 32'h00812783;
mem['h0713] = 32'h00878793;
mem['h0714] = 32'h00078593;
mem['h0715] = 32'h00040513;
mem['h0716] = 32'hEC9FF0EF;
mem['h0717] = 32'h00C12783;
mem['h0718] = 32'h0087A423;
mem['h0719] = 32'h00400513;
mem['h071A] = 32'hE31FF0EF;
mem['h071B] = 32'h00050793;
mem['h071C] = 32'h00078413;
mem['h071D] = 32'h00812783;
mem['h071E] = 32'h00C78793;
mem['h071F] = 32'h00078593;
mem['h0720] = 32'h00040513;
mem['h0721] = 32'hEC1FF0EF;
mem['h0722] = 32'h00C12783;
mem['h0723] = 32'h0087A623;
mem['h0724] = 32'h00400513;
mem['h0725] = 32'hE05FF0EF;
mem['h0726] = 32'h00050793;
mem['h0727] = 32'h00078413;
mem['h0728] = 32'h00812783;
mem['h0729] = 32'h01078793;
mem['h072A] = 32'h00078593;
mem['h072B] = 32'h00040513;
mem['h072C] = 32'hEB9FF0EF;
mem['h072D] = 32'h00C12783;
mem['h072E] = 32'h0087A823;
mem['h072F] = 32'h00400513;
mem['h0730] = 32'hDD9FF0EF;
mem['h0731] = 32'h00050793;
mem['h0732] = 32'h00078413;
mem['h0733] = 32'h00812783;
mem['h0734] = 32'h01478793;
mem['h0735] = 32'h00078593;
mem['h0736] = 32'h00040513;
mem['h0737] = 32'hEB1FF0EF;
mem['h0738] = 32'h00C12783;
mem['h0739] = 32'h0087AA23;
mem['h073A] = 32'h00400513;
mem['h073B] = 32'hDADFF0EF;
mem['h073C] = 32'h00050793;
mem['h073D] = 32'h00078413;
mem['h073E] = 32'h00812783;
mem['h073F] = 32'h01878793;
mem['h0740] = 32'h00078593;
mem['h0741] = 32'h00040513;
mem['h0742] = 32'hEA9FF0EF;
mem['h0743] = 32'h00C12783;
mem['h0744] = 32'h0087AC23;
mem['h0745] = 32'h00000013;
mem['h0746] = 32'h01C12083;
mem['h0747] = 32'h01812403;
mem['h0748] = 32'h02010113;
mem['h0749] = 32'h00008067;
mem['h074A] = 32'hFF010113;
mem['h074B] = 32'h00A12623;
mem['h074C] = 32'h00B12423;
mem['h074D] = 32'h00C12783;
mem['h074E] = 32'h00812703;
mem['h074F] = 32'h00E7A023;
mem['h0750] = 32'h00000013;
mem['h0751] = 32'h01010113;
mem['h0752] = 32'h00008067;
mem['h0753] = 32'hFF010113;
mem['h0754] = 32'h00A12623;
mem['h0755] = 32'h00B12423;
mem['h0756] = 32'h00C12783;
mem['h0757] = 32'h00812703;
mem['h0758] = 32'h00E7A023;
mem['h0759] = 32'h00000013;
mem['h075A] = 32'h01010113;
mem['h075B] = 32'h00008067;
mem['h075C] = 32'hFF010113;
mem['h075D] = 32'h00A12623;
mem['h075E] = 32'h00B12423;
mem['h075F] = 32'h00C12783;
mem['h0760] = 32'h00812703;
mem['h0761] = 32'h00E7A023;
mem['h0762] = 32'h00000013;
mem['h0763] = 32'h01010113;
mem['h0764] = 32'h00008067;
mem['h0765] = 32'hFF010113;
mem['h0766] = 32'h00A12623;
mem['h0767] = 32'h00B12423;
mem['h0768] = 32'h00C12783;
mem['h0769] = 32'h00812703;
mem['h076A] = 32'h00E7A023;
mem['h076B] = 32'h00000013;
mem['h076C] = 32'h01010113;
mem['h076D] = 32'h00008067;
mem['h076E] = 32'hFF010113;
mem['h076F] = 32'h00A12623;
mem['h0770] = 32'h00B12423;
mem['h0771] = 32'h00C12783;
mem['h0772] = 32'h00812703;
mem['h0773] = 32'h00E7A023;
mem['h0774] = 32'h00000013;
mem['h0775] = 32'h01010113;
mem['h0776] = 32'h00008067;
mem['h0777] = 32'hFF010113;
mem['h0778] = 32'h00A12623;
mem['h0779] = 32'h00B12423;
mem['h077A] = 32'h00C12783;
mem['h077B] = 32'h00812703;
mem['h077C] = 32'h00E7A023;
mem['h077D] = 32'h00000013;
mem['h077E] = 32'h01010113;
mem['h077F] = 32'h00008067;
mem['h0780] = 32'hFF010113;
mem['h0781] = 32'h00A12623;
mem['h0782] = 32'h00B12423;
mem['h0783] = 32'h00C12783;
mem['h0784] = 32'h00812703;
mem['h0785] = 32'h00E7A023;
mem['h0786] = 32'h00000013;
mem['h0787] = 32'h01010113;
mem['h0788] = 32'h00008067;
mem['h0789] = 32'hFE010113;
mem['h078A] = 32'h00112E23;
mem['h078B] = 32'h00812C23;
mem['h078C] = 32'h00A12623;
mem['h078D] = 32'h00B12423;
mem['h078E] = 32'h00400513;
mem['h078F] = 32'hC5DFF0EF;
mem['h0790] = 32'h00050793;
mem['h0791] = 32'h00078413;
mem['h0792] = 32'h00812583;
mem['h0793] = 32'h00040513;
mem['h0794] = 32'hED9FF0EF;
mem['h0795] = 32'h00C12783;
mem['h0796] = 32'h0087A023;
mem['h0797] = 32'h00400513;
mem['h0798] = 32'hC39FF0EF;
mem['h0799] = 32'h00050793;
mem['h079A] = 32'h00078413;
mem['h079B] = 32'h00812783;
mem['h079C] = 32'h00478793;
mem['h079D] = 32'h00078593;
mem['h079E] = 32'h00040513;
mem['h079F] = 32'hED1FF0EF;
mem['h07A0] = 32'h00C12783;
mem['h07A1] = 32'h0087A223;
mem['h07A2] = 32'h00400513;
mem['h07A3] = 32'hC0DFF0EF;
mem['h07A4] = 32'h00050793;
mem['h07A5] = 32'h00078413;
mem['h07A6] = 32'h00812783;
mem['h07A7] = 32'h00878793;
mem['h07A8] = 32'h00078593;
mem['h07A9] = 32'h00040513;
mem['h07AA] = 32'hEC9FF0EF;
mem['h07AB] = 32'h00C12783;
mem['h07AC] = 32'h0087A423;
mem['h07AD] = 32'h00400513;
mem['h07AE] = 32'hBE1FF0EF;
mem['h07AF] = 32'h00050793;
mem['h07B0] = 32'h00078413;
mem['h07B1] = 32'h00812783;
mem['h07B2] = 32'h00C78793;
mem['h07B3] = 32'h00078593;
mem['h07B4] = 32'h00040513;
mem['h07B5] = 32'hEC1FF0EF;
mem['h07B6] = 32'h00C12783;
mem['h07B7] = 32'h0087A623;
mem['h07B8] = 32'h00400513;
mem['h07B9] = 32'hBB5FF0EF;
mem['h07BA] = 32'h00050793;
mem['h07BB] = 32'h00078413;
mem['h07BC] = 32'h00812783;
mem['h07BD] = 32'h01078793;
mem['h07BE] = 32'h00078593;
mem['h07BF] = 32'h00040513;
mem['h07C0] = 32'hEB9FF0EF;
mem['h07C1] = 32'h00C12783;
mem['h07C2] = 32'h0087A823;
mem['h07C3] = 32'h00400513;
mem['h07C4] = 32'hB89FF0EF;
mem['h07C5] = 32'h00050793;
mem['h07C6] = 32'h00078413;
mem['h07C7] = 32'h00812783;
mem['h07C8] = 32'h01478793;
mem['h07C9] = 32'h00078593;
mem['h07CA] = 32'h00040513;
mem['h07CB] = 32'hEB1FF0EF;
mem['h07CC] = 32'h00C12783;
mem['h07CD] = 32'h0087AA23;
mem['h07CE] = 32'h00400513;
mem['h07CF] = 32'hB5DFF0EF;
mem['h07D0] = 32'h00050793;
mem['h07D1] = 32'h00078413;
mem['h07D2] = 32'h00812783;
mem['h07D3] = 32'h01878793;
mem['h07D4] = 32'h00078593;
mem['h07D5] = 32'h00040513;
mem['h07D6] = 32'hEA9FF0EF;
mem['h07D7] = 32'h00C12783;
mem['h07D8] = 32'h0087AC23;
mem['h07D9] = 32'h00000013;
mem['h07DA] = 32'h01C12083;
mem['h07DB] = 32'h01812403;
mem['h07DC] = 32'h02010113;
mem['h07DD] = 32'h00008067;
mem['h07DE] = 32'hFE010113;
mem['h07DF] = 32'h00112E23;
mem['h07E0] = 32'h00812C23;
mem['h07E1] = 32'h00A12623;
mem['h07E2] = 32'h00B12423;
mem['h07E3] = 32'h01C00513;
mem['h07E4] = 32'hB09FF0EF;
mem['h07E5] = 32'h00050793;
mem['h07E6] = 32'h00078413;
mem['h07E7] = 32'h00812583;
mem['h07E8] = 32'h00040513;
mem['h07E9] = 32'hC31FF0EF;
mem['h07EA] = 32'h00C12783;
mem['h07EB] = 32'h0087A023;
mem['h07EC] = 32'h01C00513;
mem['h07ED] = 32'hAE5FF0EF;
mem['h07EE] = 32'h00050793;
mem['h07EF] = 32'h00078413;
mem['h07F0] = 32'h00812783;
mem['h07F1] = 32'h01C78793;
mem['h07F2] = 32'h00078593;
mem['h07F3] = 32'h00040513;
mem['h07F4] = 32'hE55FF0EF;
mem['h07F5] = 32'h00C12783;
mem['h07F6] = 32'h0087A223;
mem['h07F7] = 32'h00000013;
mem['h07F8] = 32'h01C12083;
mem['h07F9] = 32'h01812403;
mem['h07FA] = 32'h02010113;
mem['h07FB] = 32'h00008067;
mem['h07FC] = 32'hFF010113;
mem['h07FD] = 32'h00A12623;
mem['h07FE] = 32'h00B12423;
mem['h07FF] = 32'h00C12783;
mem['h0800] = 32'h00812703;
mem['h0801] = 32'h00E7A023;
mem['h0802] = 32'h00000013;
mem['h0803] = 32'h01010113;
mem['h0804] = 32'h00008067;
mem['h0805] = 32'hFF010113;
mem['h0806] = 32'h00A12623;
mem['h0807] = 32'h00B12423;
mem['h0808] = 32'h00C12783;
mem['h0809] = 32'h00812703;
mem['h080A] = 32'h00E7A023;
mem['h080B] = 32'h00000013;
mem['h080C] = 32'h01010113;
mem['h080D] = 32'h00008067;
mem['h080E] = 32'hFF010113;
mem['h080F] = 32'h00A12623;
mem['h0810] = 32'h00B12423;
mem['h0811] = 32'h00C12783;
mem['h0812] = 32'h00812703;
mem['h0813] = 32'h00E7A023;
mem['h0814] = 32'h00000013;
mem['h0815] = 32'h01010113;
mem['h0816] = 32'h00008067;
mem['h0817] = 32'hFF010113;
mem['h0818] = 32'h00A12623;
mem['h0819] = 32'h00B12423;
mem['h081A] = 32'h00C12783;
mem['h081B] = 32'h00812703;
mem['h081C] = 32'h00E7A023;
mem['h081D] = 32'h00000013;
mem['h081E] = 32'h01010113;
mem['h081F] = 32'h00008067;
mem['h0820] = 32'hFE010113;
mem['h0821] = 32'h00112E23;
mem['h0822] = 32'h00812C23;
mem['h0823] = 32'h00A12623;
mem['h0824] = 32'h00B12423;
mem['h0825] = 32'h00400513;
mem['h0826] = 32'hA01FF0EF;
mem['h0827] = 32'h00050793;
mem['h0828] = 32'h00078413;
mem['h0829] = 32'h00812583;
mem['h082A] = 32'h00040513;
mem['h082B] = 32'hF45FF0EF;
mem['h082C] = 32'h00C12783;
mem['h082D] = 32'h0087A023;
mem['h082E] = 32'h00400513;
mem['h082F] = 32'h9DDFF0EF;
mem['h0830] = 32'h00050793;
mem['h0831] = 32'h00078413;
mem['h0832] = 32'h00812783;
mem['h0833] = 32'h00478793;
mem['h0834] = 32'h00078593;
mem['h0835] = 32'h00040513;
mem['h0836] = 32'hF3DFF0EF;
mem['h0837] = 32'h00C12783;
mem['h0838] = 32'h0087A223;
mem['h0839] = 32'h00400513;
mem['h083A] = 32'h9B1FF0EF;
mem['h083B] = 32'h00050793;
mem['h083C] = 32'h00078413;
mem['h083D] = 32'h00812783;
mem['h083E] = 32'h00878793;
mem['h083F] = 32'h00078593;
mem['h0840] = 32'h00040513;
mem['h0841] = 32'hF35FF0EF;
mem['h0842] = 32'h00C12783;
mem['h0843] = 32'h0087A423;
mem['h0844] = 32'h00400513;
mem['h0845] = 32'h985FF0EF;
mem['h0846] = 32'h00050793;
mem['h0847] = 32'h00078413;
mem['h0848] = 32'h00812783;
mem['h0849] = 32'h00C78793;
mem['h084A] = 32'h00078593;
mem['h084B] = 32'h00040513;
mem['h084C] = 32'hF2DFF0EF;
mem['h084D] = 32'h00C12783;
mem['h084E] = 32'h0087A623;
mem['h084F] = 32'h00000013;
mem['h0850] = 32'h01C12083;
mem['h0851] = 32'h01812403;
mem['h0852] = 32'h02010113;
mem['h0853] = 32'h00008067;
mem['h0854] = 32'hFF010113;
mem['h0855] = 32'h00A12623;
mem['h0856] = 32'h00B12423;
mem['h0857] = 32'h00C12783;
mem['h0858] = 32'h00812703;
mem['h0859] = 32'h00E7A023;
mem['h085A] = 32'h00000013;
mem['h085B] = 32'h01010113;
mem['h085C] = 32'h00008067;
mem['h085D] = 32'hFF010113;
mem['h085E] = 32'h00A12623;
mem['h085F] = 32'h00C12783;
mem['h0860] = 32'h0007A783;
mem['h0861] = 32'h0007A783;
mem['h0862] = 32'h0017F793;
mem['h0863] = 32'h0FF7F793;
mem['h0864] = 32'h00078513;
mem['h0865] = 32'h01010113;
mem['h0866] = 32'h00008067;
mem['h0867] = 32'hFF010113;
mem['h0868] = 32'h00A12623;
mem['h0869] = 32'h00B12423;
mem['h086A] = 32'h00C12783;
mem['h086B] = 32'h0007A783;
mem['h086C] = 32'h00812703;
mem['h086D] = 32'h00177713;
mem['h086E] = 32'h0FF77713;
mem['h086F] = 32'h00177713;
mem['h0870] = 32'h00871713;
mem['h0871] = 32'h0007A683;
mem['h0872] = 32'hEFF6F693;
mem['h0873] = 32'h00E6E733;
mem['h0874] = 32'h00E7A023;
mem['h0875] = 32'h00000013;
mem['h0876] = 32'h01010113;
mem['h0877] = 32'h00008067;
mem['h0878] = 32'hFF010113;
mem['h0879] = 32'h00A12623;
mem['h087A] = 32'h00B12423;
mem['h087B] = 32'h00C12783;
mem['h087C] = 32'h0007A783;
mem['h087D] = 32'h00812703;
mem['h087E] = 32'h00177713;
mem['h087F] = 32'h0FF77713;
mem['h0880] = 32'h00177713;
mem['h0881] = 32'h00971713;
mem['h0882] = 32'h0007A683;
mem['h0883] = 32'hDFF6F693;
mem['h0884] = 32'h00E6E733;
mem['h0885] = 32'h00E7A023;
mem['h0886] = 32'h00000013;
mem['h0887] = 32'h01010113;
mem['h0888] = 32'h00008067;
mem['h0889] = 32'hFF010113;
mem['h088A] = 32'h00A12623;
mem['h088B] = 32'h00B12423;
mem['h088C] = 32'h00C12783;
mem['h088D] = 32'h00812703;
mem['h088E] = 32'h00E7A023;
mem['h088F] = 32'h00000013;
mem['h0890] = 32'h01010113;
mem['h0891] = 32'h00008067;
mem['h0892] = 32'hFE010113;
mem['h0893] = 32'h00112E23;
mem['h0894] = 32'h00812C23;
mem['h0895] = 32'h00A12623;
mem['h0896] = 32'h00B12423;
mem['h0897] = 32'h00400513;
mem['h0898] = 32'h839FF0EF;
mem['h0899] = 32'h00050793;
mem['h089A] = 32'h00078413;
mem['h089B] = 32'h00812583;
mem['h089C] = 32'h00040513;
mem['h089D] = 32'hFB1FF0EF;
mem['h089E] = 32'h00C12783;
mem['h089F] = 32'h0087A023;
mem['h08A0] = 32'h00000013;
mem['h08A1] = 32'h01C12083;
mem['h08A2] = 32'h01812403;
mem['h08A3] = 32'h02010113;
mem['h08A4] = 32'h00008067;
mem['h08A5] = 32'hFF010113;
mem['h08A6] = 32'h00A12623;
mem['h08A7] = 32'h00B12423;
mem['h08A8] = 32'h00C12783;
mem['h08A9] = 32'h00812703;
mem['h08AA] = 32'h00E7A023;
mem['h08AB] = 32'h00000013;
mem['h08AC] = 32'h01010113;
mem['h08AD] = 32'h00008067;
mem['h08AE] = 32'hFE010113;
mem['h08AF] = 32'h00112E23;
mem['h08B0] = 32'h00812C23;
mem['h08B1] = 32'h00A12623;
mem['h08B2] = 32'h00B12423;
mem['h08B3] = 32'h00400513;
mem['h08B4] = 32'hFC8FF0EF;
mem['h08B5] = 32'h00050793;
mem['h08B6] = 32'h00078413;
mem['h08B7] = 32'h00812583;
mem['h08B8] = 32'h00040513;
mem['h08B9] = 32'hFB1FF0EF;
mem['h08BA] = 32'h00C12783;
mem['h08BB] = 32'h0087A023;
mem['h08BC] = 32'h00000013;
mem['h08BD] = 32'h01C12083;
mem['h08BE] = 32'h01812403;
mem['h08BF] = 32'h02010113;
mem['h08C0] = 32'h00008067;
mem['h08C1] = 32'hFF010113;
mem['h08C2] = 32'h00A12623;
mem['h08C3] = 32'h00B12423;
mem['h08C4] = 32'h00C12783;
mem['h08C5] = 32'h00812703;
mem['h08C6] = 32'h00E7A023;
mem['h08C7] = 32'h00000013;
mem['h08C8] = 32'h01010113;
mem['h08C9] = 32'h00008067;
mem['h08CA] = 32'hFD010113;
mem['h08CB] = 32'h02112623;
mem['h08CC] = 32'h02812423;
mem['h08CD] = 32'h00A12623;
mem['h08CE] = 32'h00B12423;
mem['h08CF] = 32'h00800513;
mem['h08D0] = 32'hF58FF0EF;
mem['h08D1] = 32'h00050793;
mem['h08D2] = 32'h00078413;
mem['h08D3] = 32'h00812583;
mem['h08D4] = 32'h00040513;
mem['h08D5] = 32'hC25FF0EF;
mem['h08D6] = 32'h00C12783;
mem['h08D7] = 32'h0087A023;
mem['h08D8] = 32'h01000513;
mem['h08D9] = 32'hF34FF0EF;
mem['h08DA] = 32'h00050793;
mem['h08DB] = 32'h00078413;
mem['h08DC] = 32'h00812783;
mem['h08DD] = 32'h03878793;
mem['h08DE] = 32'h00078593;
mem['h08DF] = 32'h00040513;
mem['h08E0] = 32'hD01FF0EF;
mem['h08E1] = 32'h00C12783;
mem['h08E2] = 32'h0087A223;
mem['h08E3] = 32'h00400513;
mem['h08E4] = 32'hF08FF0EF;
mem['h08E5] = 32'h00050793;
mem['h08E6] = 32'h00078413;
mem['h08E7] = 32'h00812783;
mem['h08E8] = 32'h04878793;
mem['h08E9] = 32'h00078593;
mem['h08EA] = 32'h00040513;
mem['h08EB] = 32'hDA5FF0EF;
mem['h08EC] = 32'h00C12783;
mem['h08ED] = 32'h0087A423;
mem['h08EE] = 32'h00012E23;
mem['h08EF] = 32'h0540006F;
mem['h08F0] = 32'h00400513;
mem['h08F1] = 32'hED4FF0EF;
mem['h08F2] = 32'h00050793;
mem['h08F3] = 32'h00078413;
mem['h08F4] = 32'h01C12783;
mem['h08F5] = 32'h01378793;
mem['h08F6] = 32'h00279793;
mem['h08F7] = 32'h00812703;
mem['h08F8] = 32'h00F707B3;
mem['h08F9] = 32'h00078593;
mem['h08FA] = 32'h00040513;
mem['h08FB] = 32'hE5DFF0EF;
mem['h08FC] = 32'h00C12703;
mem['h08FD] = 32'h01C12783;
mem['h08FE] = 32'h00279793;
mem['h08FF] = 32'h00F707B3;
mem['h0900] = 32'h0087A623;
mem['h0901] = 32'h01C12783;
mem['h0902] = 32'h00178793;
mem['h0903] = 32'h00F12E23;
mem['h0904] = 32'h01C12703;
mem['h0905] = 32'h00300793;
mem['h0906] = 32'hFAE7D4E3;
mem['h0907] = 32'h00400513;
mem['h0908] = 32'hE78FF0EF;
mem['h0909] = 32'h00050793;
mem['h090A] = 32'h00078413;
mem['h090B] = 32'h00812783;
mem['h090C] = 32'h05C78793;
mem['h090D] = 32'h00078593;
mem['h090E] = 32'h00040513;
mem['h090F] = 32'hE7DFF0EF;
mem['h0910] = 32'h00C12783;
mem['h0911] = 32'h0087AE23;
mem['h0912] = 32'h00400513;
mem['h0913] = 32'hE4CFF0EF;
mem['h0914] = 32'h00050793;
mem['h0915] = 32'h00078413;
mem['h0916] = 32'h00812783;
mem['h0917] = 32'h06078793;
mem['h0918] = 32'h00078593;
mem['h0919] = 32'h00040513;
mem['h091A] = 32'hE9DFF0EF;
mem['h091B] = 32'h00C12783;
mem['h091C] = 32'h0287A023;
mem['h091D] = 32'h00000013;
mem['h091E] = 32'h02C12083;
mem['h091F] = 32'h02812403;
mem['h0920] = 32'h03010113;
mem['h0921] = 32'h00008067;
mem['h0922] = 32'hFB010113;
mem['h0923] = 32'h04112623;
mem['h0924] = 32'h04812423;
mem['h0925] = 32'h02400513;
mem['h0926] = 32'hE00FF0EF;
mem['h0927] = 32'h00050793;
mem['h0928] = 32'h00078413;
mem['h0929] = 32'h200005B7;
mem['h092A] = 32'h00040513;
mem['h092B] = 32'hE7DFF0EF;
mem['h092C] = 32'h02812C23;
mem['h092D] = 32'h03812783;
mem['h092E] = 32'h0087A783;
mem['h092F] = 32'h00100593;
mem['h0930] = 32'h00078513;
mem['h0931] = 32'hD1DFF0EF;
mem['h0932] = 32'h03812783;
mem['h0933] = 32'h0087A403;
mem['h0934] = 32'h03812783;
mem['h0935] = 32'h0087A783;
mem['h0936] = 32'h00078513;
mem['h0937] = 32'hC99FF0EF;
mem['h0938] = 32'h00050793;
mem['h0939] = 32'h00078593;
mem['h093A] = 32'h00040513;
mem['h093B] = 32'hCB1FF0EF;
mem['h093C] = 32'h000027B7;
mem['h093D] = 32'h74878793;
mem['h093E] = 32'h0007A603;
mem['h093F] = 32'h0047A683;
mem['h0940] = 32'h0087A703;
mem['h0941] = 32'h00C12423;
mem['h0942] = 32'h00D12623;
mem['h0943] = 32'h00E12823;
mem['h0944] = 32'h00C7D703;
mem['h0945] = 32'h00E11A23;
mem['h0946] = 32'h00E7C783;
mem['h0947] = 32'h00F10B23;
mem['h0948] = 32'h00810793;
mem['h0949] = 32'h02F12E23;
mem['h094A] = 32'h0200006F;
mem['h094B] = 32'h03C12783;
mem['h094C] = 32'h00178713;
mem['h094D] = 32'h02E12E23;
mem['h094E] = 32'h0007C783;
mem['h094F] = 32'h00078593;
mem['h0950] = 32'h03812503;
mem['h0951] = 32'hBA1FD0EF;
mem['h0952] = 32'h03C12783;
mem['h0953] = 32'h0007C783;
mem['h0954] = 32'hFC079EE3;
mem['h0955] = 32'h00000793;
mem['h0956] = 32'h00078513;
mem['h0957] = 32'h04C12083;
mem['h0958] = 32'h04812403;
mem['h0959] = 32'h05010113;
mem['h095A] = 32'h00008067;
mem['h095B] = 32'h00050613;
mem['h095C] = 32'h00000513;
mem['h095D] = 32'h0015F693;
mem['h095E] = 32'h00068463;
mem['h095F] = 32'h00C50533;
mem['h0960] = 32'h0015D593;
mem['h0961] = 32'h00161613;
mem['h0962] = 32'hFE0596E3;
mem['h0963] = 32'h00008067;
mem['h0964] = 32'h06054063;
mem['h0965] = 32'h0605C663;
mem['h0966] = 32'h00058613;
mem['h0967] = 32'h00050593;
mem['h0968] = 32'hFFF00513;
mem['h0969] = 32'h02060C63;
mem['h096A] = 32'h00100693;
mem['h096B] = 32'h00B67A63;
mem['h096C] = 32'h00C05863;
mem['h096D] = 32'h00161613;
mem['h096E] = 32'h00169693;
mem['h096F] = 32'hFEB66AE3;
mem['h0970] = 32'h00000513;
mem['h0971] = 32'h00C5E663;
mem['h0972] = 32'h40C585B3;
mem['h0973] = 32'h00D56533;
mem['h0974] = 32'h0016D693;
mem['h0975] = 32'h00165613;
mem['h0976] = 32'hFE0696E3;
mem['h0977] = 32'h00008067;
mem['h0978] = 32'h00008293;
mem['h0979] = 32'hFB5FF0EF;
mem['h097A] = 32'h00058513;
mem['h097B] = 32'h00028067;
mem['h097C] = 32'h40A00533;
mem['h097D] = 32'h00B04863;
mem['h097E] = 32'h40B005B3;
mem['h097F] = 32'hF9DFF06F;
mem['h0980] = 32'h40B005B3;
mem['h0981] = 32'h00008293;
mem['h0982] = 32'hF91FF0EF;
mem['h0983] = 32'h40A00533;
mem['h0984] = 32'h00028067;
mem['h0985] = 32'h00008293;
mem['h0986] = 32'h0005CA63;
mem['h0987] = 32'h00054C63;
mem['h0988] = 32'hF79FF0EF;
mem['h0989] = 32'h00058513;
mem['h098A] = 32'h00028067;
mem['h098B] = 32'h40B005B3;
mem['h098C] = 32'hFE0558E3;
mem['h098D] = 32'h40A00533;
mem['h098E] = 32'hF61FF0EF;
mem['h098F] = 32'h40B00533;
mem['h0990] = 32'h00028067;
mem['h0991] = 32'h33323130;
mem['h0992] = 32'h37363534;
mem['h0993] = 32'h42413938;
mem['h0994] = 32'h46454443;
mem['h0995] = 32'h00000000;
mem['h0996] = 32'h7320694D;
mem['h0997] = 32'h46206F6D;
mem['h0998] = 32'h20414750;
mem['h0999] = 32'h616A6172;
mem['h099A] = 32'h00000000;
mem['h099B] = 32'h530A0A0D;
mem['h099C] = 32'h6D616C65;
mem['h099D] = 32'h75646520;
mem['h099E] = 32'h20434F53;
mem['h099F] = 32'h6B636148;
mem['h09A0] = 32'h21737265;
mem['h09A1] = 32'h00000A0D;
mem['h09A2] = 32'h20797254;
mem['h09A3] = 32'h73657567;
mem['h09A4] = 32'h676E6973;
mem['h09A5] = 32'h74203320;
mem['h09A6] = 32'h73656D69;
mem['h09A7] = 32'h61687720;
mem['h09A8] = 32'h27492074;
mem['h09A9] = 32'h6874206D;
mem['h09AA] = 32'h696B6E69;
mem['h09AB] = 32'h202C676E;
mem['h09AC] = 32'h6E656874;
mem['h09AD] = 32'h65727020;
mem['h09AE] = 32'h3C207373;
mem['h09AF] = 32'h45544E45;
mem['h09B0] = 32'h0D2E3E52;
mem['h09B1] = 32'h0000000A;
mem['h09B2] = 32'h090A0A0D;
mem['h09B3] = 32'h20756F59;
mem['h09B4] = 32'h65746E65;
mem['h09B5] = 32'h3A646572;
mem['h09B6] = 32'h00000020;
mem['h09B7] = 32'h7C090A0D;
mem['h09B8] = 32'h756F5920;
mem['h09B9] = 32'h74696820;
mem['h09BA] = 32'h21746920;
mem['h09BB] = 32'h292D3A20;
mem['h09BC] = 32'h00000A0D;
mem['h09BD] = 32'h7C090A0D;
mem['h09BE] = 32'h726F5320;
mem['h09BF] = 32'h202C7972;
mem['h09C0] = 32'h20756F79;
mem['h09C1] = 32'h7373696D;
mem['h09C2] = 32'h69206465;
mem['h09C3] = 32'h00002E74;
mem['h09C4] = 32'h7C090A0D;
mem['h09C5] = 32'h2E2E2E20;
mem['h09C6] = 32'h20797254;
mem['h09C7] = 32'h69616761;
mem['h09C8] = 32'h43202E6E;
mem['h09C9] = 32'h69646572;
mem['h09CA] = 32'h656C2074;
mem['h09CB] = 32'h203A7466;
mem['h09CC] = 32'h00000000;
mem['h09CD] = 32'h0A0A0A0D;
mem['h09CE] = 32'h00000000;
mem['h09CF] = 32'h4F440A0D;
mem['h09D0] = 32'h0D21454E;
mem['h09D1] = 32'h0000000A;
mem['h09D2] = 32'h6C6C6548;
mem['h09D3] = 32'h6F77206F;
mem['h09D4] = 32'h21646C72;
mem['h09D5] = 32'h00000A0D;
