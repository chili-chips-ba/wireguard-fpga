mem['h0000] = 32'h00001517;
mem['h0001] = 32'hBB850513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h00418593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h0E0000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'hFE010113;
mem['h001D] = 32'h00A12623;
mem['h001E] = 32'h0001A783;
mem['h001F] = 32'h00078713;
mem['h0020] = 32'h100007B7;
mem['h0021] = 32'h00078793;
mem['h0022] = 32'h00F707B3;
mem['h0023] = 32'h00F12E23;
mem['h0024] = 32'h0001A703;
mem['h0025] = 32'h00C12783;
mem['h0026] = 32'h00F70733;
mem['h0027] = 32'h00E1A023;
mem['h0028] = 32'h0001A703;
mem['h0029] = 32'h000017B7;
mem['h002A] = 32'h80078793;
mem['h002B] = 32'h00E7D463;
mem['h002C] = 32'h00100073;
mem['h002D] = 32'h01C12783;
mem['h002E] = 32'h00078513;
mem['h002F] = 32'h02010113;
mem['h0030] = 32'h00008067;
mem['h0031] = 32'hFD010113;
mem['h0032] = 32'h02112623;
mem['h0033] = 32'h00A12623;
mem['h0034] = 32'h00C12783;
mem['h0035] = 32'h00078513;
mem['h0036] = 32'hF99FF0EF;
mem['h0037] = 32'h00A12E23;
mem['h0038] = 32'h01C12783;
mem['h0039] = 32'h00078513;
mem['h003A] = 32'h02C12083;
mem['h003B] = 32'h03010113;
mem['h003C] = 32'h00008067;
mem['h003D] = 32'hFF010113;
mem['h003E] = 32'h00A12623;
mem['h003F] = 32'h00000013;
mem['h0040] = 32'h01010113;
mem['h0041] = 32'h00008067;
mem['h0042] = 32'hFE010113;
mem['h0043] = 32'h00A12623;
mem['h0044] = 32'h00012E23;
mem['h0045] = 32'h0100006F;
mem['h0046] = 32'h01C12783;
mem['h0047] = 32'h00178793;
mem['h0048] = 32'h00F12E23;
mem['h0049] = 32'h01C12783;
mem['h004A] = 32'h00C12703;
mem['h004B] = 32'h00E7B7B3;
mem['h004C] = 32'h0FF7F793;
mem['h004D] = 32'hFE0792E3;
mem['h004E] = 32'h00000013;
mem['h004F] = 32'h00000013;
mem['h0050] = 32'h02010113;
mem['h0051] = 32'h00008067;
mem['h0052] = 32'hFE010113;
mem['h0053] = 32'h00112E23;
mem['h0054] = 32'h00812C23;
mem['h0055] = 32'h02400513;
mem['h0056] = 32'hF6DFF0EF;
mem['h0057] = 32'h00050793;
mem['h0058] = 32'h00078413;
mem['h0059] = 32'h200005B7;
mem['h005A] = 32'h00040513;
mem['h005B] = 32'h0ED000EF;
mem['h005C] = 32'h00812623;
mem['h005D] = 32'h00C12783;
mem['h005E] = 32'h0087A783;
mem['h005F] = 32'h00100593;
mem['h0060] = 32'h00078513;
mem['h0061] = 32'h78C000EF;
mem['h0062] = 32'h00C12783;
mem['h0063] = 32'h0087A403;
mem['h0064] = 32'h00C12783;
mem['h0065] = 32'h0087A783;
mem['h0066] = 32'h00078513;
mem['h0067] = 32'h708000EF;
mem['h0068] = 32'h00050793;
mem['h0069] = 32'h00078593;
mem['h006A] = 32'h00040513;
mem['h006B] = 32'h720000EF;
mem['h006C] = 32'h000F47B7;
mem['h006D] = 32'h24078513;
mem['h006E] = 32'hF51FF0EF;
mem['h006F] = 32'h00C12783;
mem['h0070] = 32'h0087A783;
mem['h0071] = 32'h00000593;
mem['h0072] = 32'h00078513;
mem['h0073] = 32'h744000EF;
mem['h0074] = 32'h00C12783;
mem['h0075] = 32'h0087A403;
mem['h0076] = 32'h00C12783;
mem['h0077] = 32'h0087A783;
mem['h0078] = 32'h00078513;
mem['h0079] = 32'h6C0000EF;
mem['h007A] = 32'h00050793;
mem['h007B] = 32'h00078593;
mem['h007C] = 32'h00040513;
mem['h007D] = 32'h6D8000EF;
mem['h007E] = 32'h000F47B7;
mem['h007F] = 32'h24078513;
mem['h0080] = 32'hF09FF0EF;
mem['h0081] = 32'hF71FF06F;
mem['h0082] = 32'hFF010113;
mem['h0083] = 32'h00A12623;
mem['h0084] = 32'h00B12423;
mem['h0085] = 32'h00C12783;
mem['h0086] = 32'h00812703;
mem['h0087] = 32'h00E7A023;
mem['h0088] = 32'h00000013;
mem['h0089] = 32'h01010113;
mem['h008A] = 32'h00008067;
mem['h008B] = 32'hFF010113;
mem['h008C] = 32'h00A12623;
mem['h008D] = 32'h00B12423;
mem['h008E] = 32'h00C12783;
mem['h008F] = 32'h00812703;
mem['h0090] = 32'h00E7A023;
mem['h0091] = 32'h00000013;
mem['h0092] = 32'h01010113;
mem['h0093] = 32'h00008067;
mem['h0094] = 32'hFF010113;
mem['h0095] = 32'h00A12623;
mem['h0096] = 32'h00B12423;
mem['h0097] = 32'h00C12783;
mem['h0098] = 32'h00812703;
mem['h0099] = 32'h00E7A023;
mem['h009A] = 32'h00000013;
mem['h009B] = 32'h01010113;
mem['h009C] = 32'h00008067;
mem['h009D] = 32'hFF010113;
mem['h009E] = 32'h00A12623;
mem['h009F] = 32'h00B12423;
mem['h00A0] = 32'h00C12783;
mem['h00A1] = 32'h00812703;
mem['h00A2] = 32'h00E7A023;
mem['h00A3] = 32'h00000013;
mem['h00A4] = 32'h01010113;
mem['h00A5] = 32'h00008067;
mem['h00A6] = 32'hFF010113;
mem['h00A7] = 32'h00A12623;
mem['h00A8] = 32'h00B12423;
mem['h00A9] = 32'h00C12783;
mem['h00AA] = 32'h00812703;
mem['h00AB] = 32'h00E7A023;
mem['h00AC] = 32'h00000013;
mem['h00AD] = 32'h01010113;
mem['h00AE] = 32'h00008067;
mem['h00AF] = 32'hFF010113;
mem['h00B0] = 32'h00A12623;
mem['h00B1] = 32'h00B12423;
mem['h00B2] = 32'h00C12783;
mem['h00B3] = 32'h00812703;
mem['h00B4] = 32'h00E7A023;
mem['h00B5] = 32'h00000013;
mem['h00B6] = 32'h01010113;
mem['h00B7] = 32'h00008067;
mem['h00B8] = 32'hFF010113;
mem['h00B9] = 32'h00A12623;
mem['h00BA] = 32'h00B12423;
mem['h00BB] = 32'h00C12783;
mem['h00BC] = 32'h00812703;
mem['h00BD] = 32'h00E7A023;
mem['h00BE] = 32'h00000013;
mem['h00BF] = 32'h01010113;
mem['h00C0] = 32'h00008067;
mem['h00C1] = 32'hFE010113;
mem['h00C2] = 32'h00112E23;
mem['h00C3] = 32'h00812C23;
mem['h00C4] = 32'h00A12623;
mem['h00C5] = 32'h00B12423;
mem['h00C6] = 32'h00400513;
mem['h00C7] = 32'hDA9FF0EF;
mem['h00C8] = 32'h00050793;
mem['h00C9] = 32'h00078413;
mem['h00CA] = 32'h00812583;
mem['h00CB] = 32'h00040513;
mem['h00CC] = 32'hED9FF0EF;
mem['h00CD] = 32'h00C12783;
mem['h00CE] = 32'h0087A023;
mem['h00CF] = 32'h00400513;
mem['h00D0] = 32'hD85FF0EF;
mem['h00D1] = 32'h00050793;
mem['h00D2] = 32'h00078413;
mem['h00D3] = 32'h00812783;
mem['h00D4] = 32'h00478793;
mem['h00D5] = 32'h00078593;
mem['h00D6] = 32'h00040513;
mem['h00D7] = 32'hED1FF0EF;
mem['h00D8] = 32'h00C12783;
mem['h00D9] = 32'h0087A223;
mem['h00DA] = 32'h00400513;
mem['h00DB] = 32'hD59FF0EF;
mem['h00DC] = 32'h00050793;
mem['h00DD] = 32'h00078413;
mem['h00DE] = 32'h00812783;
mem['h00DF] = 32'h00878793;
mem['h00E0] = 32'h00078593;
mem['h00E1] = 32'h00040513;
mem['h00E2] = 32'hEC9FF0EF;
mem['h00E3] = 32'h00C12783;
mem['h00E4] = 32'h0087A423;
mem['h00E5] = 32'h00400513;
mem['h00E6] = 32'hD2DFF0EF;
mem['h00E7] = 32'h00050793;
mem['h00E8] = 32'h00078413;
mem['h00E9] = 32'h00812783;
mem['h00EA] = 32'h00C78793;
mem['h00EB] = 32'h00078593;
mem['h00EC] = 32'h00040513;
mem['h00ED] = 32'hEC1FF0EF;
mem['h00EE] = 32'h00C12783;
mem['h00EF] = 32'h0087A623;
mem['h00F0] = 32'h00400513;
mem['h00F1] = 32'hD01FF0EF;
mem['h00F2] = 32'h00050793;
mem['h00F3] = 32'h00078413;
mem['h00F4] = 32'h00812783;
mem['h00F5] = 32'h01078793;
mem['h00F6] = 32'h00078593;
mem['h00F7] = 32'h00040513;
mem['h00F8] = 32'hEB9FF0EF;
mem['h00F9] = 32'h00C12783;
mem['h00FA] = 32'h0087A823;
mem['h00FB] = 32'h00400513;
mem['h00FC] = 32'hCD5FF0EF;
mem['h00FD] = 32'h00050793;
mem['h00FE] = 32'h00078413;
mem['h00FF] = 32'h00812783;
mem['h0100] = 32'h01478793;
mem['h0101] = 32'h00078593;
mem['h0102] = 32'h00040513;
mem['h0103] = 32'hEB1FF0EF;
mem['h0104] = 32'h00C12783;
mem['h0105] = 32'h0087AA23;
mem['h0106] = 32'h00400513;
mem['h0107] = 32'hCA9FF0EF;
mem['h0108] = 32'h00050793;
mem['h0109] = 32'h00078413;
mem['h010A] = 32'h00812783;
mem['h010B] = 32'h01878793;
mem['h010C] = 32'h00078593;
mem['h010D] = 32'h00040513;
mem['h010E] = 32'hEA9FF0EF;
mem['h010F] = 32'h00C12783;
mem['h0110] = 32'h0087AC23;
mem['h0111] = 32'h00000013;
mem['h0112] = 32'h01C12083;
mem['h0113] = 32'h01812403;
mem['h0114] = 32'h02010113;
mem['h0115] = 32'h00008067;
mem['h0116] = 32'hFF010113;
mem['h0117] = 32'h00A12623;
mem['h0118] = 32'h00B12423;
mem['h0119] = 32'h00C12783;
mem['h011A] = 32'h00812703;
mem['h011B] = 32'h00E7A023;
mem['h011C] = 32'h00000013;
mem['h011D] = 32'h01010113;
mem['h011E] = 32'h00008067;
mem['h011F] = 32'hFF010113;
mem['h0120] = 32'h00A12623;
mem['h0121] = 32'h00B12423;
mem['h0122] = 32'h00C12783;
mem['h0123] = 32'h00812703;
mem['h0124] = 32'h00E7A023;
mem['h0125] = 32'h00000013;
mem['h0126] = 32'h01010113;
mem['h0127] = 32'h00008067;
mem['h0128] = 32'hFF010113;
mem['h0129] = 32'h00A12623;
mem['h012A] = 32'h00B12423;
mem['h012B] = 32'h00C12783;
mem['h012C] = 32'h00812703;
mem['h012D] = 32'h00E7A023;
mem['h012E] = 32'h00000013;
mem['h012F] = 32'h01010113;
mem['h0130] = 32'h00008067;
mem['h0131] = 32'hFF010113;
mem['h0132] = 32'h00A12623;
mem['h0133] = 32'h00B12423;
mem['h0134] = 32'h00C12783;
mem['h0135] = 32'h00812703;
mem['h0136] = 32'h00E7A023;
mem['h0137] = 32'h00000013;
mem['h0138] = 32'h01010113;
mem['h0139] = 32'h00008067;
mem['h013A] = 32'hFF010113;
mem['h013B] = 32'h00A12623;
mem['h013C] = 32'h00B12423;
mem['h013D] = 32'h00C12783;
mem['h013E] = 32'h00812703;
mem['h013F] = 32'h00E7A023;
mem['h0140] = 32'h00000013;
mem['h0141] = 32'h01010113;
mem['h0142] = 32'h00008067;
mem['h0143] = 32'hFF010113;
mem['h0144] = 32'h00A12623;
mem['h0145] = 32'h00B12423;
mem['h0146] = 32'h00C12783;
mem['h0147] = 32'h00812703;
mem['h0148] = 32'h00E7A023;
mem['h0149] = 32'h00000013;
mem['h014A] = 32'h01010113;
mem['h014B] = 32'h00008067;
mem['h014C] = 32'hFF010113;
mem['h014D] = 32'h00A12623;
mem['h014E] = 32'h00B12423;
mem['h014F] = 32'h00C12783;
mem['h0150] = 32'h00812703;
mem['h0151] = 32'h00E7A023;
mem['h0152] = 32'h00000013;
mem['h0153] = 32'h01010113;
mem['h0154] = 32'h00008067;
mem['h0155] = 32'hFE010113;
mem['h0156] = 32'h00112E23;
mem['h0157] = 32'h00812C23;
mem['h0158] = 32'h00A12623;
mem['h0159] = 32'h00B12423;
mem['h015A] = 32'h00400513;
mem['h015B] = 32'hB59FF0EF;
mem['h015C] = 32'h00050793;
mem['h015D] = 32'h00078413;
mem['h015E] = 32'h00812583;
mem['h015F] = 32'h00040513;
mem['h0160] = 32'hED9FF0EF;
mem['h0161] = 32'h00C12783;
mem['h0162] = 32'h0087A023;
mem['h0163] = 32'h00400513;
mem['h0164] = 32'hB35FF0EF;
mem['h0165] = 32'h00050793;
mem['h0166] = 32'h00078413;
mem['h0167] = 32'h00812783;
mem['h0168] = 32'h00478793;
mem['h0169] = 32'h00078593;
mem['h016A] = 32'h00040513;
mem['h016B] = 32'hED1FF0EF;
mem['h016C] = 32'h00C12783;
mem['h016D] = 32'h0087A223;
mem['h016E] = 32'h00400513;
mem['h016F] = 32'hB09FF0EF;
mem['h0170] = 32'h00050793;
mem['h0171] = 32'h00078413;
mem['h0172] = 32'h00812783;
mem['h0173] = 32'h00878793;
mem['h0174] = 32'h00078593;
mem['h0175] = 32'h00040513;
mem['h0176] = 32'hEC9FF0EF;
mem['h0177] = 32'h00C12783;
mem['h0178] = 32'h0087A423;
mem['h0179] = 32'h00400513;
mem['h017A] = 32'hADDFF0EF;
mem['h017B] = 32'h00050793;
mem['h017C] = 32'h00078413;
mem['h017D] = 32'h00812783;
mem['h017E] = 32'h00C78793;
mem['h017F] = 32'h00078593;
mem['h0180] = 32'h00040513;
mem['h0181] = 32'hEC1FF0EF;
mem['h0182] = 32'h00C12783;
mem['h0183] = 32'h0087A623;
mem['h0184] = 32'h00400513;
mem['h0185] = 32'hAB1FF0EF;
mem['h0186] = 32'h00050793;
mem['h0187] = 32'h00078413;
mem['h0188] = 32'h00812783;
mem['h0189] = 32'h01078793;
mem['h018A] = 32'h00078593;
mem['h018B] = 32'h00040513;
mem['h018C] = 32'hEB9FF0EF;
mem['h018D] = 32'h00C12783;
mem['h018E] = 32'h0087A823;
mem['h018F] = 32'h00400513;
mem['h0190] = 32'hA85FF0EF;
mem['h0191] = 32'h00050793;
mem['h0192] = 32'h00078413;
mem['h0193] = 32'h00812783;
mem['h0194] = 32'h01478793;
mem['h0195] = 32'h00078593;
mem['h0196] = 32'h00040513;
mem['h0197] = 32'hEB1FF0EF;
mem['h0198] = 32'h00C12783;
mem['h0199] = 32'h0087AA23;
mem['h019A] = 32'h00400513;
mem['h019B] = 32'hA59FF0EF;
mem['h019C] = 32'h00050793;
mem['h019D] = 32'h00078413;
mem['h019E] = 32'h00812783;
mem['h019F] = 32'h01878793;
mem['h01A0] = 32'h00078593;
mem['h01A1] = 32'h00040513;
mem['h01A2] = 32'hEA9FF0EF;
mem['h01A3] = 32'h00C12783;
mem['h01A4] = 32'h0087AC23;
mem['h01A5] = 32'h00000013;
mem['h01A6] = 32'h01C12083;
mem['h01A7] = 32'h01812403;
mem['h01A8] = 32'h02010113;
mem['h01A9] = 32'h00008067;
mem['h01AA] = 32'hFE010113;
mem['h01AB] = 32'h00112E23;
mem['h01AC] = 32'h00812C23;
mem['h01AD] = 32'h00A12623;
mem['h01AE] = 32'h00B12423;
mem['h01AF] = 32'h01C00513;
mem['h01B0] = 32'hA05FF0EF;
mem['h01B1] = 32'h00050793;
mem['h01B2] = 32'h00078413;
mem['h01B3] = 32'h00812583;
mem['h01B4] = 32'h00040513;
mem['h01B5] = 32'hC31FF0EF;
mem['h01B6] = 32'h00C12783;
mem['h01B7] = 32'h0087A023;
mem['h01B8] = 32'h01C00513;
mem['h01B9] = 32'h9E1FF0EF;
mem['h01BA] = 32'h00050793;
mem['h01BB] = 32'h00078413;
mem['h01BC] = 32'h00812783;
mem['h01BD] = 32'h01C78793;
mem['h01BE] = 32'h00078593;
mem['h01BF] = 32'h00040513;
mem['h01C0] = 32'hE55FF0EF;
mem['h01C1] = 32'h00C12783;
mem['h01C2] = 32'h0087A223;
mem['h01C3] = 32'h00000013;
mem['h01C4] = 32'h01C12083;
mem['h01C5] = 32'h01812403;
mem['h01C6] = 32'h02010113;
mem['h01C7] = 32'h00008067;
mem['h01C8] = 32'hFF010113;
mem['h01C9] = 32'h00A12623;
mem['h01CA] = 32'h00B12423;
mem['h01CB] = 32'h00C12783;
mem['h01CC] = 32'h00812703;
mem['h01CD] = 32'h00E7A023;
mem['h01CE] = 32'h00000013;
mem['h01CF] = 32'h01010113;
mem['h01D0] = 32'h00008067;
mem['h01D1] = 32'hFF010113;
mem['h01D2] = 32'h00A12623;
mem['h01D3] = 32'h00B12423;
mem['h01D4] = 32'h00C12783;
mem['h01D5] = 32'h00812703;
mem['h01D6] = 32'h00E7A023;
mem['h01D7] = 32'h00000013;
mem['h01D8] = 32'h01010113;
mem['h01D9] = 32'h00008067;
mem['h01DA] = 32'hFF010113;
mem['h01DB] = 32'h00A12623;
mem['h01DC] = 32'h00B12423;
mem['h01DD] = 32'h00C12783;
mem['h01DE] = 32'h00812703;
mem['h01DF] = 32'h00E7A023;
mem['h01E0] = 32'h00000013;
mem['h01E1] = 32'h01010113;
mem['h01E2] = 32'h00008067;
mem['h01E3] = 32'hFF010113;
mem['h01E4] = 32'h00A12623;
mem['h01E5] = 32'h00B12423;
mem['h01E6] = 32'h00C12783;
mem['h01E7] = 32'h00812703;
mem['h01E8] = 32'h00E7A023;
mem['h01E9] = 32'h00000013;
mem['h01EA] = 32'h01010113;
mem['h01EB] = 32'h00008067;
mem['h01EC] = 32'hFE010113;
mem['h01ED] = 32'h00112E23;
mem['h01EE] = 32'h00812C23;
mem['h01EF] = 32'h00A12623;
mem['h01F0] = 32'h00B12423;
mem['h01F1] = 32'h00400513;
mem['h01F2] = 32'h8FDFF0EF;
mem['h01F3] = 32'h00050793;
mem['h01F4] = 32'h00078413;
mem['h01F5] = 32'h00812583;
mem['h01F6] = 32'h00040513;
mem['h01F7] = 32'hF45FF0EF;
mem['h01F8] = 32'h00C12783;
mem['h01F9] = 32'h0087A023;
mem['h01FA] = 32'h00400513;
mem['h01FB] = 32'h8D9FF0EF;
mem['h01FC] = 32'h00050793;
mem['h01FD] = 32'h00078413;
mem['h01FE] = 32'h00812783;
mem['h01FF] = 32'h00478793;
mem['h0200] = 32'h00078593;
mem['h0201] = 32'h00040513;
mem['h0202] = 32'hF3DFF0EF;
mem['h0203] = 32'h00C12783;
mem['h0204] = 32'h0087A223;
mem['h0205] = 32'h00400513;
mem['h0206] = 32'h8ADFF0EF;
mem['h0207] = 32'h00050793;
mem['h0208] = 32'h00078413;
mem['h0209] = 32'h00812783;
mem['h020A] = 32'h00878793;
mem['h020B] = 32'h00078593;
mem['h020C] = 32'h00040513;
mem['h020D] = 32'hF35FF0EF;
mem['h020E] = 32'h00C12783;
mem['h020F] = 32'h0087A423;
mem['h0210] = 32'h00400513;
mem['h0211] = 32'h881FF0EF;
mem['h0212] = 32'h00050793;
mem['h0213] = 32'h00078413;
mem['h0214] = 32'h00812783;
mem['h0215] = 32'h00C78793;
mem['h0216] = 32'h00078593;
mem['h0217] = 32'h00040513;
mem['h0218] = 32'hF2DFF0EF;
mem['h0219] = 32'h00C12783;
mem['h021A] = 32'h0087A623;
mem['h021B] = 32'h00000013;
mem['h021C] = 32'h01C12083;
mem['h021D] = 32'h01812403;
mem['h021E] = 32'h02010113;
mem['h021F] = 32'h00008067;
mem['h0220] = 32'hFF010113;
mem['h0221] = 32'h00A12623;
mem['h0222] = 32'h00B12423;
mem['h0223] = 32'h00C12783;
mem['h0224] = 32'h00812703;
mem['h0225] = 32'h00E7A023;
mem['h0226] = 32'h00000013;
mem['h0227] = 32'h01010113;
mem['h0228] = 32'h00008067;
mem['h0229] = 32'hFF010113;
mem['h022A] = 32'h00A12623;
mem['h022B] = 32'h00C12783;
mem['h022C] = 32'h0007A783;
mem['h022D] = 32'h0007A783;
mem['h022E] = 32'h0017F793;
mem['h022F] = 32'h0FF7F793;
mem['h0230] = 32'h00078513;
mem['h0231] = 32'h01010113;
mem['h0232] = 32'h00008067;
mem['h0233] = 32'hFF010113;
mem['h0234] = 32'h00A12623;
mem['h0235] = 32'h00B12423;
mem['h0236] = 32'h00C12783;
mem['h0237] = 32'h0007A783;
mem['h0238] = 32'h00812703;
mem['h0239] = 32'h00177713;
mem['h023A] = 32'h0FF77713;
mem['h023B] = 32'h00177713;
mem['h023C] = 32'h00871713;
mem['h023D] = 32'h0007A683;
mem['h023E] = 32'hEFF6F693;
mem['h023F] = 32'h00E6E733;
mem['h0240] = 32'h00E7A023;
mem['h0241] = 32'h00000013;
mem['h0242] = 32'h01010113;
mem['h0243] = 32'h00008067;
mem['h0244] = 32'hFF010113;
mem['h0245] = 32'h00A12623;
mem['h0246] = 32'h00B12423;
mem['h0247] = 32'h00C12783;
mem['h0248] = 32'h0007A783;
mem['h0249] = 32'h00812703;
mem['h024A] = 32'h00177713;
mem['h024B] = 32'h0FF77713;
mem['h024C] = 32'h00177713;
mem['h024D] = 32'h00971713;
mem['h024E] = 32'h0007A683;
mem['h024F] = 32'hDFF6F693;
mem['h0250] = 32'h00E6E733;
mem['h0251] = 32'h00E7A023;
mem['h0252] = 32'h00000013;
mem['h0253] = 32'h01010113;
mem['h0254] = 32'h00008067;
mem['h0255] = 32'hFF010113;
mem['h0256] = 32'h00A12623;
mem['h0257] = 32'h00B12423;
mem['h0258] = 32'h00C12783;
mem['h0259] = 32'h00812703;
mem['h025A] = 32'h00E7A023;
mem['h025B] = 32'h00000013;
mem['h025C] = 32'h01010113;
mem['h025D] = 32'h00008067;
mem['h025E] = 32'hFE010113;
mem['h025F] = 32'h00112E23;
mem['h0260] = 32'h00812C23;
mem['h0261] = 32'h00A12623;
mem['h0262] = 32'h00B12423;
mem['h0263] = 32'h00400513;
mem['h0264] = 32'hF34FF0EF;
mem['h0265] = 32'h00050793;
mem['h0266] = 32'h00078413;
mem['h0267] = 32'h00812583;
mem['h0268] = 32'h00040513;
mem['h0269] = 32'hFB1FF0EF;
mem['h026A] = 32'h00C12783;
mem['h026B] = 32'h0087A023;
mem['h026C] = 32'h00000013;
mem['h026D] = 32'h01C12083;
mem['h026E] = 32'h01812403;
mem['h026F] = 32'h02010113;
mem['h0270] = 32'h00008067;
mem['h0271] = 32'hFF010113;
mem['h0272] = 32'h00A12623;
mem['h0273] = 32'h00B12423;
mem['h0274] = 32'h00C12783;
mem['h0275] = 32'h00812703;
mem['h0276] = 32'h00E7A023;
mem['h0277] = 32'h00000013;
mem['h0278] = 32'h01010113;
mem['h0279] = 32'h00008067;
mem['h027A] = 32'hFE010113;
mem['h027B] = 32'h00112E23;
mem['h027C] = 32'h00812C23;
mem['h027D] = 32'h00A12623;
mem['h027E] = 32'h00B12423;
mem['h027F] = 32'h00400513;
mem['h0280] = 32'hEC4FF0EF;
mem['h0281] = 32'h00050793;
mem['h0282] = 32'h00078413;
mem['h0283] = 32'h00812583;
mem['h0284] = 32'h00040513;
mem['h0285] = 32'hFB1FF0EF;
mem['h0286] = 32'h00C12783;
mem['h0287] = 32'h0087A023;
mem['h0288] = 32'h00000013;
mem['h0289] = 32'h01C12083;
mem['h028A] = 32'h01812403;
mem['h028B] = 32'h02010113;
mem['h028C] = 32'h00008067;
mem['h028D] = 32'hFF010113;
mem['h028E] = 32'h00A12623;
mem['h028F] = 32'h00B12423;
mem['h0290] = 32'h00C12783;
mem['h0291] = 32'h00812703;
mem['h0292] = 32'h00E7A023;
mem['h0293] = 32'h00000013;
mem['h0294] = 32'h01010113;
mem['h0295] = 32'h00008067;
mem['h0296] = 32'hFD010113;
mem['h0297] = 32'h02112623;
mem['h0298] = 32'h02812423;
mem['h0299] = 32'h00A12623;
mem['h029A] = 32'h00B12423;
mem['h029B] = 32'h00800513;
mem['h029C] = 32'hE54FF0EF;
mem['h029D] = 32'h00050793;
mem['h029E] = 32'h00078413;
mem['h029F] = 32'h00812583;
mem['h02A0] = 32'h00040513;
mem['h02A1] = 32'hC25FF0EF;
mem['h02A2] = 32'h00C12783;
mem['h02A3] = 32'h0087A023;
mem['h02A4] = 32'h01000513;
mem['h02A5] = 32'hE30FF0EF;
mem['h02A6] = 32'h00050793;
mem['h02A7] = 32'h00078413;
mem['h02A8] = 32'h00812783;
mem['h02A9] = 32'h03878793;
mem['h02AA] = 32'h00078593;
mem['h02AB] = 32'h00040513;
mem['h02AC] = 32'hD01FF0EF;
mem['h02AD] = 32'h00C12783;
mem['h02AE] = 32'h0087A223;
mem['h02AF] = 32'h00400513;
mem['h02B0] = 32'hE04FF0EF;
mem['h02B1] = 32'h00050793;
mem['h02B2] = 32'h00078413;
mem['h02B3] = 32'h00812783;
mem['h02B4] = 32'h04878793;
mem['h02B5] = 32'h00078593;
mem['h02B6] = 32'h00040513;
mem['h02B7] = 32'hDA5FF0EF;
mem['h02B8] = 32'h00C12783;
mem['h02B9] = 32'h0087A423;
mem['h02BA] = 32'h00012E23;
mem['h02BB] = 32'h0540006F;
mem['h02BC] = 32'h00400513;
mem['h02BD] = 32'hDD0FF0EF;
mem['h02BE] = 32'h00050793;
mem['h02BF] = 32'h00078413;
mem['h02C0] = 32'h01C12783;
mem['h02C1] = 32'h01378793;
mem['h02C2] = 32'h00279793;
mem['h02C3] = 32'h00812703;
mem['h02C4] = 32'h00F707B3;
mem['h02C5] = 32'h00078593;
mem['h02C6] = 32'h00040513;
mem['h02C7] = 32'hE5DFF0EF;
mem['h02C8] = 32'h00C12703;
mem['h02C9] = 32'h01C12783;
mem['h02CA] = 32'h00279793;
mem['h02CB] = 32'h00F707B3;
mem['h02CC] = 32'h0087A623;
mem['h02CD] = 32'h01C12783;
mem['h02CE] = 32'h00178793;
mem['h02CF] = 32'h00F12E23;
mem['h02D0] = 32'h01C12703;
mem['h02D1] = 32'h00300793;
mem['h02D2] = 32'hFAE7D4E3;
mem['h02D3] = 32'h00400513;
mem['h02D4] = 32'hD74FF0EF;
mem['h02D5] = 32'h00050793;
mem['h02D6] = 32'h00078413;
mem['h02D7] = 32'h00812783;
mem['h02D8] = 32'h05C78793;
mem['h02D9] = 32'h00078593;
mem['h02DA] = 32'h00040513;
mem['h02DB] = 32'hE7DFF0EF;
mem['h02DC] = 32'h00C12783;
mem['h02DD] = 32'h0087AE23;
mem['h02DE] = 32'h00400513;
mem['h02DF] = 32'hD48FF0EF;
mem['h02E0] = 32'h00050793;
mem['h02E1] = 32'h00078413;
mem['h02E2] = 32'h00812783;
mem['h02E3] = 32'h06078793;
mem['h02E4] = 32'h00078593;
mem['h02E5] = 32'h00040513;
mem['h02E6] = 32'hE9DFF0EF;
mem['h02E7] = 32'h00C12783;
mem['h02E8] = 32'h0287A023;
mem['h02E9] = 32'h00000013;
mem['h02EA] = 32'h02C12083;
mem['h02EB] = 32'h02812403;
mem['h02EC] = 32'h03010113;
mem['h02ED] = 32'h00008067;
