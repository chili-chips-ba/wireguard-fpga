-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity chacha20_state_to_bytes_0CLK_d3fba2d7 is
port(
 x : in chacha20_state;
 return_output : out uint8_t_array_64_t);
end chacha20_state_to_bytes_0CLK_d3fba2d7;
architecture arch of chacha20_state_to_bytes_0CLK_d3fba2d7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065]
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
signal FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;

function CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned) return uint8_t_array_64_t is
 
  variable base : uint8_t_array_64_t; 
  variable return_output : uint8_t_array_64_t;
begin
      base.data(0) := ref_toks_0;
      base.data(1) := ref_toks_1;
      base.data(2) := ref_toks_2;
      base.data(3) := ref_toks_3;
      base.data(4) := ref_toks_4;
      base.data(5) := ref_toks_5;
      base.data(6) := ref_toks_6;
      base.data(7) := ref_toks_7;
      base.data(8) := ref_toks_8;
      base.data(9) := ref_toks_9;
      base.data(10) := ref_toks_10;
      base.data(11) := ref_toks_11;
      base.data(12) := ref_toks_12;
      base.data(13) := ref_toks_13;
      base.data(14) := ref_toks_14;
      base.data(15) := ref_toks_15;
      base.data(16) := ref_toks_16;
      base.data(17) := ref_toks_17;
      base.data(18) := ref_toks_18;
      base.data(19) := ref_toks_19;
      base.data(20) := ref_toks_20;
      base.data(21) := ref_toks_21;
      base.data(22) := ref_toks_22;
      base.data(23) := ref_toks_23;
      base.data(24) := ref_toks_24;
      base.data(25) := ref_toks_25;
      base.data(26) := ref_toks_26;
      base.data(27) := ref_toks_27;
      base.data(28) := ref_toks_28;
      base.data(29) := ref_toks_29;
      base.data(30) := ref_toks_30;
      base.data(31) := ref_toks_31;
      base.data(32) := ref_toks_32;
      base.data(33) := ref_toks_33;
      base.data(34) := ref_toks_34;
      base.data(35) := ref_toks_35;
      base.data(36) := ref_toks_36;
      base.data(37) := ref_toks_37;
      base.data(38) := ref_toks_38;
      base.data(39) := ref_toks_39;
      base.data(40) := ref_toks_40;
      base.data(41) := ref_toks_41;
      base.data(42) := ref_toks_42;
      base.data(43) := ref_toks_43;
      base.data(44) := ref_toks_44;
      base.data(45) := ref_toks_45;
      base.data(46) := ref_toks_46;
      base.data(47) := ref_toks_47;
      base.data(48) := ref_toks_48;
      base.data(49) := ref_toks_49;
      base.data(50) := ref_toks_50;
      base.data(51) := ref_toks_51;
      base.data(52) := ref_toks_52;
      base.data(53) := ref_toks_53;
      base.data(54) := ref_toks_54;
      base.data(55) := ref_toks_55;
      base.data(56) := ref_toks_56;
      base.data(57) := ref_toks_57;
      base.data(58) := ref_toks_58;
      base.data(59) := ref_toks_59;
      base.data(60) := ref_toks_60;
      base.data(61) := ref_toks_61;
      base.data(62) := ref_toks_62;
      base.data(63) := ref_toks_63;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);

-- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : 0 clocks latency
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065 : entity work.uint32_t_to_bytes_0CLK_a5a1cd4e port map (
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x,
FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 x,
 -- All submodule outputs
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output,
 FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : uint8_t_array_64_t;
 variable VAR_x : chacha20_state;
 variable VAR_rv : uint8_t_array_64_t;
 variable VAR_pos : unsigned(6 downto 0);
 variable VAR_field_pos : unsigned(6 downto 0);
 variable VAR_state_dim_0 : unsigned(4 downto 0);
 variable VAR_state_elem_bytes : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output : uint8_t_array_4_t;
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef_chacha20_state_bytes_t_h_l25_c12_c130_return_output : uint8_t_array_64_t;
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_x := x;

     -- Submodule level 0
     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(13);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(15);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(7);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(9);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(10);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(11);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(4);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(14);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(8);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(6);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(5);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d[chacha20_state_bytes_t_h_l17_c57_8a88] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output := VAR_x.state(12);

     -- Submodule level 1
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_CONST_REF_RD_uint32_t_chacha20_state_state_0_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_CONST_REF_RD_uint32_t_chacha20_state_state_10_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_CONST_REF_RD_uint32_t_chacha20_state_state_11_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_CONST_REF_RD_uint32_t_chacha20_state_state_12_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_CONST_REF_RD_uint32_t_chacha20_state_state_13_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_CONST_REF_RD_uint32_t_chacha20_state_state_14_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_CONST_REF_RD_uint32_t_chacha20_state_state_15_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_CONST_REF_RD_uint32_t_chacha20_state_state_1_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_CONST_REF_RD_uint32_t_chacha20_state_state_2_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_CONST_REF_RD_uint32_t_chacha20_state_state_3_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_CONST_REF_RD_uint32_t_chacha20_state_state_4_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_CONST_REF_RD_uint32_t_chacha20_state_state_5_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_CONST_REF_RD_uint32_t_chacha20_state_state_6_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_CONST_REF_RD_uint32_t_chacha20_state_state_7_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_CONST_REF_RD_uint32_t_chacha20_state_state_8_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_CONST_REF_RD_uint32_t_chacha20_state_state_9_d41d_chacha20_state_bytes_t_h_l17_c57_8a88_return_output;
     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes[chacha20_state_bytes_t_h_l17_c39_3065] LATENCY=0
     -- Inputs
     FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x <= VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_x;
     -- Outputs
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output := FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output;

     -- Submodule level 2
     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(3);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(1);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(2);

     -- FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d[chacha20_state_bytes_t_h_l20_c20_2229] LATENCY=0
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output := VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_uint32_t_to_bytes_chacha20_state_bytes_t_h_l17_c39_3065_return_output.data(0);

     -- Submodule level 3
     -- CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef[chacha20_state_bytes_t_h_l25_c12_c130] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef_chacha20_state_bytes_t_h_l25_c12_c130_return_output := CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef(
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_0_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_1_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_2_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_3_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_4_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_5_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_6_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_7_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_8_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_9_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_10_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_11_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_12_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_13_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_14_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_0_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_1_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_2_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output,
     VAR_FOR_chacha20_state_bytes_t_h_l16_c1_f5a8_ITER_15_FOR_chacha20_state_bytes_t_h_l18_c2_e5e8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_array_4_t_data_3_d41d_chacha20_state_bytes_t_h_l20_c20_2229_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_64_t_uint8_t_array_64_t_f9ef_chacha20_state_bytes_t_h_l25_c12_c130_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
