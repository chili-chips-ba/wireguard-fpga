-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 7
entity axis512_to_axis128_array_0CLK_4b8d8b28 is
port(
 axis : in axis512_t;
 return_output : out axis512_to_axis128_array_t);
end axis512_to_axis128_array_0CLK_4b8d8b28;
architecture arch of axis512_to_axis128_array_0CLK_4b8d8b28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT[axis_h_l329_c36_f263]
signal FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND[axis_h_l330_c35_b026]
signal FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT[axis_h_l329_c36_f263]
signal FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND[axis_h_l330_c35_b026]
signal FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT[axis_h_l329_c36_f263]
signal FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND[axis_h_l330_c35_b026]
signal FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
signal FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);

function CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned;
 ref_toks_113 : unsigned;
 ref_toks_114 : unsigned;
 ref_toks_115 : unsigned;
 ref_toks_116 : unsigned;
 ref_toks_117 : unsigned;
 ref_toks_118 : unsigned;
 ref_toks_119 : unsigned;
 ref_toks_120 : unsigned;
 ref_toks_121 : unsigned;
 ref_toks_122 : unsigned;
 ref_toks_123 : unsigned;
 ref_toks_124 : unsigned;
 ref_toks_125 : unsigned;
 ref_toks_126 : unsigned;
 ref_toks_127 : unsigned;
 ref_toks_128 : unsigned;
 ref_toks_129 : unsigned;
 ref_toks_130 : unsigned;
 ref_toks_131 : unsigned;
 ref_toks_132 : unsigned;
 ref_toks_133 : unsigned;
 ref_toks_134 : unsigned;
 ref_toks_135 : unsigned) return axis512_to_axis128_array_t is
 
  variable base : axis512_to_axis128_array_t; 
  variable return_output : axis512_to_axis128_array_t;
begin
      base.axis_chunks(0).valid := ref_toks_0;
      base.axis_chunks(0).data.tdata(0) := ref_toks_1;
      base.axis_chunks(0).data.tkeep(0) := ref_toks_2;
      base.axis_chunks(0).data.tdata(1) := ref_toks_3;
      base.axis_chunks(0).data.tkeep(1) := ref_toks_4;
      base.axis_chunks(0).data.tdata(2) := ref_toks_5;
      base.axis_chunks(0).data.tkeep(2) := ref_toks_6;
      base.axis_chunks(0).data.tdata(3) := ref_toks_7;
      base.axis_chunks(0).data.tkeep(3) := ref_toks_8;
      base.axis_chunks(0).data.tdata(4) := ref_toks_9;
      base.axis_chunks(0).data.tkeep(4) := ref_toks_10;
      base.axis_chunks(0).data.tdata(5) := ref_toks_11;
      base.axis_chunks(0).data.tkeep(5) := ref_toks_12;
      base.axis_chunks(0).data.tdata(6) := ref_toks_13;
      base.axis_chunks(0).data.tkeep(6) := ref_toks_14;
      base.axis_chunks(0).data.tdata(7) := ref_toks_15;
      base.axis_chunks(0).data.tkeep(7) := ref_toks_16;
      base.axis_chunks(0).data.tdata(8) := ref_toks_17;
      base.axis_chunks(0).data.tkeep(8) := ref_toks_18;
      base.axis_chunks(0).data.tdata(9) := ref_toks_19;
      base.axis_chunks(0).data.tkeep(9) := ref_toks_20;
      base.axis_chunks(0).data.tdata(10) := ref_toks_21;
      base.axis_chunks(0).data.tkeep(10) := ref_toks_22;
      base.axis_chunks(0).data.tdata(11) := ref_toks_23;
      base.axis_chunks(0).data.tkeep(11) := ref_toks_24;
      base.axis_chunks(0).data.tdata(12) := ref_toks_25;
      base.axis_chunks(0).data.tkeep(12) := ref_toks_26;
      base.axis_chunks(0).data.tdata(13) := ref_toks_27;
      base.axis_chunks(0).data.tkeep(13) := ref_toks_28;
      base.axis_chunks(0).data.tdata(14) := ref_toks_29;
      base.axis_chunks(0).data.tkeep(14) := ref_toks_30;
      base.axis_chunks(0).data.tdata(15) := ref_toks_31;
      base.axis_chunks(0).data.tkeep(15) := ref_toks_32;
      base.axis_chunks(1).valid := ref_toks_33;
      base.axis_chunks(1).data.tdata(0) := ref_toks_34;
      base.axis_chunks(1).data.tkeep(0) := ref_toks_35;
      base.axis_chunks(1).data.tdata(1) := ref_toks_36;
      base.axis_chunks(1).data.tkeep(1) := ref_toks_37;
      base.axis_chunks(1).data.tdata(2) := ref_toks_38;
      base.axis_chunks(1).data.tkeep(2) := ref_toks_39;
      base.axis_chunks(1).data.tdata(3) := ref_toks_40;
      base.axis_chunks(1).data.tkeep(3) := ref_toks_41;
      base.axis_chunks(1).data.tdata(4) := ref_toks_42;
      base.axis_chunks(1).data.tkeep(4) := ref_toks_43;
      base.axis_chunks(1).data.tdata(5) := ref_toks_44;
      base.axis_chunks(1).data.tkeep(5) := ref_toks_45;
      base.axis_chunks(1).data.tdata(6) := ref_toks_46;
      base.axis_chunks(1).data.tkeep(6) := ref_toks_47;
      base.axis_chunks(1).data.tdata(7) := ref_toks_48;
      base.axis_chunks(1).data.tkeep(7) := ref_toks_49;
      base.axis_chunks(1).data.tdata(8) := ref_toks_50;
      base.axis_chunks(1).data.tkeep(8) := ref_toks_51;
      base.axis_chunks(1).data.tdata(9) := ref_toks_52;
      base.axis_chunks(1).data.tkeep(9) := ref_toks_53;
      base.axis_chunks(1).data.tdata(10) := ref_toks_54;
      base.axis_chunks(1).data.tkeep(10) := ref_toks_55;
      base.axis_chunks(1).data.tdata(11) := ref_toks_56;
      base.axis_chunks(1).data.tkeep(11) := ref_toks_57;
      base.axis_chunks(1).data.tdata(12) := ref_toks_58;
      base.axis_chunks(1).data.tkeep(12) := ref_toks_59;
      base.axis_chunks(1).data.tdata(13) := ref_toks_60;
      base.axis_chunks(1).data.tkeep(13) := ref_toks_61;
      base.axis_chunks(1).data.tdata(14) := ref_toks_62;
      base.axis_chunks(1).data.tkeep(14) := ref_toks_63;
      base.axis_chunks(1).data.tdata(15) := ref_toks_64;
      base.axis_chunks(1).data.tkeep(15) := ref_toks_65;
      base.axis_chunks(2).valid := ref_toks_66;
      base.axis_chunks(2).data.tdata(0) := ref_toks_67;
      base.axis_chunks(2).data.tkeep(0) := ref_toks_68;
      base.axis_chunks(2).data.tdata(1) := ref_toks_69;
      base.axis_chunks(2).data.tkeep(1) := ref_toks_70;
      base.axis_chunks(2).data.tdata(2) := ref_toks_71;
      base.axis_chunks(2).data.tkeep(2) := ref_toks_72;
      base.axis_chunks(2).data.tdata(3) := ref_toks_73;
      base.axis_chunks(2).data.tkeep(3) := ref_toks_74;
      base.axis_chunks(2).data.tdata(4) := ref_toks_75;
      base.axis_chunks(2).data.tkeep(4) := ref_toks_76;
      base.axis_chunks(2).data.tdata(5) := ref_toks_77;
      base.axis_chunks(2).data.tkeep(5) := ref_toks_78;
      base.axis_chunks(2).data.tdata(6) := ref_toks_79;
      base.axis_chunks(2).data.tkeep(6) := ref_toks_80;
      base.axis_chunks(2).data.tdata(7) := ref_toks_81;
      base.axis_chunks(2).data.tkeep(7) := ref_toks_82;
      base.axis_chunks(2).data.tdata(8) := ref_toks_83;
      base.axis_chunks(2).data.tkeep(8) := ref_toks_84;
      base.axis_chunks(2).data.tdata(9) := ref_toks_85;
      base.axis_chunks(2).data.tkeep(9) := ref_toks_86;
      base.axis_chunks(2).data.tdata(10) := ref_toks_87;
      base.axis_chunks(2).data.tkeep(10) := ref_toks_88;
      base.axis_chunks(2).data.tdata(11) := ref_toks_89;
      base.axis_chunks(2).data.tkeep(11) := ref_toks_90;
      base.axis_chunks(2).data.tdata(12) := ref_toks_91;
      base.axis_chunks(2).data.tkeep(12) := ref_toks_92;
      base.axis_chunks(2).data.tdata(13) := ref_toks_93;
      base.axis_chunks(2).data.tkeep(13) := ref_toks_94;
      base.axis_chunks(2).data.tdata(14) := ref_toks_95;
      base.axis_chunks(2).data.tkeep(14) := ref_toks_96;
      base.axis_chunks(2).data.tdata(15) := ref_toks_97;
      base.axis_chunks(2).data.tkeep(15) := ref_toks_98;
      base.axis_chunks(3).valid := ref_toks_99;
      base.axis_chunks(3).data.tdata(0) := ref_toks_100;
      base.axis_chunks(3).data.tkeep(0) := ref_toks_101;
      base.axis_chunks(3).data.tdata(1) := ref_toks_102;
      base.axis_chunks(3).data.tkeep(1) := ref_toks_103;
      base.axis_chunks(3).data.tdata(2) := ref_toks_104;
      base.axis_chunks(3).data.tkeep(2) := ref_toks_105;
      base.axis_chunks(3).data.tdata(3) := ref_toks_106;
      base.axis_chunks(3).data.tkeep(3) := ref_toks_107;
      base.axis_chunks(3).data.tdata(4) := ref_toks_108;
      base.axis_chunks(3).data.tkeep(4) := ref_toks_109;
      base.axis_chunks(3).data.tdata(5) := ref_toks_110;
      base.axis_chunks(3).data.tkeep(5) := ref_toks_111;
      base.axis_chunks(3).data.tdata(6) := ref_toks_112;
      base.axis_chunks(3).data.tkeep(6) := ref_toks_113;
      base.axis_chunks(3).data.tdata(7) := ref_toks_114;
      base.axis_chunks(3).data.tkeep(7) := ref_toks_115;
      base.axis_chunks(3).data.tdata(8) := ref_toks_116;
      base.axis_chunks(3).data.tkeep(8) := ref_toks_117;
      base.axis_chunks(3).data.tdata(9) := ref_toks_118;
      base.axis_chunks(3).data.tkeep(9) := ref_toks_119;
      base.axis_chunks(3).data.tdata(10) := ref_toks_120;
      base.axis_chunks(3).data.tkeep(10) := ref_toks_121;
      base.axis_chunks(3).data.tdata(11) := ref_toks_122;
      base.axis_chunks(3).data.tkeep(11) := ref_toks_123;
      base.axis_chunks(3).data.tdata(12) := ref_toks_124;
      base.axis_chunks(3).data.tkeep(12) := ref_toks_125;
      base.axis_chunks(3).data.tdata(13) := ref_toks_126;
      base.axis_chunks(3).data.tkeep(13) := ref_toks_127;
      base.axis_chunks(3).data.tdata(14) := ref_toks_128;
      base.axis_chunks(3).data.tkeep(14) := ref_toks_129;
      base.axis_chunks(3).data.tdata(15) := ref_toks_130;
      base.axis_chunks(3).data.tkeep(15) := ref_toks_131;
      base.axis_chunks(3).data.tlast := ref_toks_132;
      base.axis_chunks(0).data.tlast := ref_toks_133;
      base.axis_chunks(1).data.tlast := ref_toks_134;
      base.axis_chunks(2).data.tlast := ref_toks_135;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr,
FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output);

-- FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left,
FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right,
FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output);

-- FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr,
FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output);

-- FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left,
FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right,
FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output);

-- FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr,
FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output);

-- FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026 : 0 clocks latency
FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left,
FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right,
FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 axis,
 -- All submodule outputs
 FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output,
 FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output,
 FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output,
 FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output,
 FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output,
 FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis512_to_axis128_array_t;
 variable VAR_axis : axis512_t;
 variable VAR_o : axis512_to_axis128_array_t;
 variable VAR_CHUNK_SIZE : unsigned(31 downto 0);
 variable VAR_c : unsigned(31 downto 0);
 variable VAR_b : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_0_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_1_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_1_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_2_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_2_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_3_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_3_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_4_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_4_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_5_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_5_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_6_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_6_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_7_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_7_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_8_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_8_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_9_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_9_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_10_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_10_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_11_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_11_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_12_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_12_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_13_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_13_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_14_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_14_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_15_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_15_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_16_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_17_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_17_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_18_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_18_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_19_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_19_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_20_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_20_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_21_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_21_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_22_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_22_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_23_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_23_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_24_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_24_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_25_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_25_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_26_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_26_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_27_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_27_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_28_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_28_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_29_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_29_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_30_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_30_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_31_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_31_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_32_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_33_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_33_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_34_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_34_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_35_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_35_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_36_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_36_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_37_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_37_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_38_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_38_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_39_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_39_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_40_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_40_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_41_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_41_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_42_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_42_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_43_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_43_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_44_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_44_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_45_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_45_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_46_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_46_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_47_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_47_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_48_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_49_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_49_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_50_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_50_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_51_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_51_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_52_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_52_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_53_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_53_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_54_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_54_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_55_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_55_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_56_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_56_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_57_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_57_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_58_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_58_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_59_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_59_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_60_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_60_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_61_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_61_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_62_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_62_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_63_d41d_axis_h_l318_c40_7cee_return_output : unsigned(7 downto 0);
 variable VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_63_d41d_axis_h_l319_c40_3735_return_output : unsigned(0 downto 0);
 variable VAR_next_chunk_is_empty : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6_axis_h_l332_c10_cc76_return_output : axis512_to_axis128_array_t;
 variable VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_0_d41d_axis_h_l315_l319_DUPLICATE_38ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_axis := axis;

     -- Submodule level 0
     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_47_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_47_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(47);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_19_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_19_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(19);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_26_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_26_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(26);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_18_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_18_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(18);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_26_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_26_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(26);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_15_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_15_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(15);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_10_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_10_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(10);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_33_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_33_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(33);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_63_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_63_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(63);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_61_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_61_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(61);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_53_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_53_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(53);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_44_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_44_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(44);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_31_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_31_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(31);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_15_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_15_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(15);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_38_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_38_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(38);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_43_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_43_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(43);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_12_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_12_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(12);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_45_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_45_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(45);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_17_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_17_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(17);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_58_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_58_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(58);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_55_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_55_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(55);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_2_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_2_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(2);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_40_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_40_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(40);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_1_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_1_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(1);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_2_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_2_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(2);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_28_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_28_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(28);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_57_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_57_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(57);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_29_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_29_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(29);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_35_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_35_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(35);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_62_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_62_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(62);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_44_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_44_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(44);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_37_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_37_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(37);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_59_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_59_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(59);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_9_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_9_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(9);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_25_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_25_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(25);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_50_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_50_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(50);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_11_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_11_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(11);

     -- CONST_REF_RD_uint1_t_axis512_t_tkeep_0_d41d_axis_h_l315_l319_DUPLICATE_38ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_0_d41d_axis_h_l315_l319_DUPLICATE_38ba_return_output := VAR_axis.tkeep(0);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_16_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_16_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(16);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_6_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_6_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(6);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_3_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_3_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(3);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_7_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_7_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(7);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_5_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_5_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(5);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_40_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_40_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(40);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_34_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_34_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(34);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_43_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_43_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(43);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_56_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_56_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(56);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_51_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_51_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(51);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_48_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_48_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(48);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_6_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_6_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(6);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_14_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_14_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(14);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_50_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_50_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(50);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_25_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_25_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(25);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_63_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_63_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(63);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_21_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_21_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(21);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_5_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_5_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(5);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_20_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_20_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(20);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_35_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_35_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(35);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_11_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_11_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(11);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_9_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_9_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(9);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_21_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_21_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(21);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_28_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_28_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(28);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_7_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_7_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(7);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_8_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_8_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(8);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_18_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_18_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(18);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_36_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_36_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(36);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_30_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_30_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(30);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_30_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_30_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(30);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_52_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_52_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(52);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_55_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_55_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(55);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_46_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_46_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(46);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_47_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_47_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(47);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_41_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_41_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(41);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_60_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_60_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(60);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_57_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_57_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(57);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_54_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_54_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(54);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_27_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_27_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(27);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_45_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_45_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(45);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_33_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_33_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(33);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_58_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_58_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(58);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_19_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_19_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(19);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_42_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_42_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(42);

     -- CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output := VAR_axis.tlast;

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_60_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_60_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(60);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_20_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_20_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(20);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_39_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_39_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(39);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_51_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_51_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(51);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_53_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_53_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(53);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_24_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_24_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(24);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_13_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_13_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(13);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_36_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_36_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(36);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_10_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_10_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(10);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_4_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_4_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(4);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_1_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_1_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(1);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_31_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_31_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(31);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_12_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_12_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(12);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_38_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_38_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(38);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_56_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_56_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(56);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_0_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_0_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(0);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_14_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_14_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(14);

     -- CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5_return_output := VAR_axis.tkeep(48);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_13_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_13_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(13);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_52_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_52_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(52);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_17_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_17_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(17);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_49_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_49_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(49);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_34_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_34_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(34);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_61_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_61_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(61);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_29_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_29_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(29);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_23_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_23_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(23);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_41_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_41_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(41);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_24_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_24_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(24);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_32_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_32_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(32);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_8_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_8_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(8);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_46_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_46_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(46);

     -- CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e_return_output := VAR_axis.tkeep(32);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_39_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_39_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(39);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_62_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_62_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(62);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_42_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_42_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(42);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_22_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_22_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(22);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_22_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_22_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(22);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_4_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_4_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(4);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_23_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_23_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(23);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_49_d41d[axis_h_l319_c40_3735] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_49_d41d_axis_h_l319_c40_3735_return_output := VAR_axis.tkeep(49);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_54_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_54_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(54);

     -- FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_37_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_37_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(37);

     -- FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_27_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_27_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(27);

     -- FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_3_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_3_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(3);

     -- CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4_return_output := VAR_axis.tkeep(16);

     -- FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_59_d41d[axis_h_l318_c40_7cee] LATENCY=0
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_59_d41d_axis_h_l318_c40_7cee_return_output := VAR_axis.tdata(59);

     -- Submodule level 1
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr := VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr := VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr := VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left := VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left := VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left := VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output;
     -- FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT[axis_h_l329_c36_f263] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr <= VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_expr;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output := FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;

     -- FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT[axis_h_l329_c36_f263] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr <= VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_expr;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output := FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;

     -- FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT[axis_h_l329_c36_f263] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr <= VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_expr;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output := FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;

     -- Submodule level 2
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right := VAR_FOR_axis_h_l327_c3_3b13_ITER_0_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right := VAR_FOR_axis_h_l327_c3_3b13_ITER_1_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right := VAR_FOR_axis_h_l327_c3_3b13_ITER_2_UNARY_OP_NOT_axis_h_l329_c36_f263_return_output;
     -- FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND[axis_h_l330_c35_b026] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left <= VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_left;
     FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right <= VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_right;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output := FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output;

     -- FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND[axis_h_l330_c35_b026] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left <= VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_left;
     FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right <= VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_right;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output := FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output;

     -- FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND[axis_h_l330_c35_b026] LATENCY=0
     -- Inputs
     FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left <= VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_left;
     FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right <= VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_right;
     -- Outputs
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output := FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output;

     -- Submodule level 3
     -- CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6[axis_h_l332_c10_cc76] LATENCY=0
     VAR_CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6_axis_h_l332_c10_cc76_return_output := CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6(
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_0_d41d_axis_h_l315_l319_DUPLICATE_38ba_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_0_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_0_d41d_axis_h_l315_l319_DUPLICATE_38ba_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_1_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_1_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_2_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_2_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_3_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_3_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_4_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_4_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_5_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_5_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_6_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_6_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_7_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_7_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_8_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_8_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_9_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_9_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_10_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_10_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_11_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_11_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_12_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_12_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_13_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_13_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_14_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_14_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_15_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_0_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_15_d41d_axis_h_l319_c40_3735_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_16_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_16_d41d_axis_h_l315_l319_DUPLICATE_74d4_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_17_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_17_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_18_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_18_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_19_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_19_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_20_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_20_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_21_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_21_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_22_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_22_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_23_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_23_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_24_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_24_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_25_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_25_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_26_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_26_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_27_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_27_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_28_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_28_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_29_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_29_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_30_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_30_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_31_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_1_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_31_d41d_axis_h_l319_c40_3735_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_32_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_32_d41d_axis_h_l315_l319_DUPLICATE_762e_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_33_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_33_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_34_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_34_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_35_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_35_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_36_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_36_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_37_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_37_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_38_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_38_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_39_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_39_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_40_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_40_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_41_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_41_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_42_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_42_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_43_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_43_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_44_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_44_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_45_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_45_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_46_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_46_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_47_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_2_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_47_d41d_axis_h_l319_c40_3735_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_0_CONST_REF_RD_uint8_t_axis512_t_tdata_48_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tkeep_48_d41d_axis_h_l315_l319_DUPLICATE_d5d5_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint8_t_axis512_t_tdata_49_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_1_CONST_REF_RD_uint1_t_axis512_t_tkeep_49_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint8_t_axis512_t_tdata_50_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_2_CONST_REF_RD_uint1_t_axis512_t_tkeep_50_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint8_t_axis512_t_tdata_51_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_3_CONST_REF_RD_uint1_t_axis512_t_tkeep_51_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint8_t_axis512_t_tdata_52_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_4_CONST_REF_RD_uint1_t_axis512_t_tkeep_52_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint8_t_axis512_t_tdata_53_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_5_CONST_REF_RD_uint1_t_axis512_t_tkeep_53_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint8_t_axis512_t_tdata_54_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_6_CONST_REF_RD_uint1_t_axis512_t_tkeep_54_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint8_t_axis512_t_tdata_55_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_7_CONST_REF_RD_uint1_t_axis512_t_tkeep_55_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint8_t_axis512_t_tdata_56_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_8_CONST_REF_RD_uint1_t_axis512_t_tkeep_56_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint8_t_axis512_t_tdata_57_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_9_CONST_REF_RD_uint1_t_axis512_t_tkeep_57_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint8_t_axis512_t_tdata_58_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_10_CONST_REF_RD_uint1_t_axis512_t_tkeep_58_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint8_t_axis512_t_tdata_59_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_11_CONST_REF_RD_uint1_t_axis512_t_tkeep_59_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint8_t_axis512_t_tdata_60_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_12_CONST_REF_RD_uint1_t_axis512_t_tkeep_60_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint8_t_axis512_t_tdata_61_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_13_CONST_REF_RD_uint1_t_axis512_t_tkeep_61_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint8_t_axis512_t_tdata_62_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_14_CONST_REF_RD_uint1_t_axis512_t_tkeep_62_d41d_axis_h_l319_c40_3735_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint8_t_axis512_t_tdata_63_d41d_axis_h_l318_c40_7cee_return_output,
     VAR_FOR_axis_h_l311_c3_887e_ITER_3_FOR_axis_h_l316_c5_ec95_ITER_15_CONST_REF_RD_uint1_t_axis512_t_tkeep_63_d41d_axis_h_l319_c40_3735_return_output,
     VAR_CONST_REF_RD_uint1_t_axis512_t_tlast_d41d_axis_h_l326_l330_DUPLICATE_850a_return_output,
     VAR_FOR_axis_h_l327_c3_3b13_ITER_0_BIN_OP_AND_axis_h_l330_c35_b026_return_output,
     VAR_FOR_axis_h_l327_c3_3b13_ITER_1_BIN_OP_AND_axis_h_l330_c35_b026_return_output,
     VAR_FOR_axis_h_l327_c3_3b13_ITER_2_BIN_OP_AND_axis_h_l330_c35_b026_return_output);

     -- Submodule level 4
     VAR_return_output := VAR_CONST_REF_RD_axis512_to_axis128_array_t_axis512_to_axis128_array_t_b4f6_axis_h_l332_c10_cc76_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
